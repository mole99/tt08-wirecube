// SPDX-FileCopyrightText: © 2024 Leo Moser <leo.moser@pm.me>
// SPDX-License-Identifier: Apache-2.0

`default_nettype none

module line_rom (
    input  logic [4:0] frame_i, // 32 frames
    input  logic [3:0] line_i,  // 12 lines
    
    output types::line_t      my_line,
    output logic [types::THRESH_BITS-1:0] my_thresh
);
    // Line
    always_comb begin
        case (line_i)
            4'd0: my_line = line_0[frame_i];
            4'd1: my_line = line_1[frame_i];
            4'd2: my_line = line_2[frame_i];
            4'd3: my_line = line_3[frame_i];
            4'd4: my_line = line_4[frame_i];
            4'd5: my_line = line_5[frame_i];
            4'd6: my_line = line_6[frame_i];
            4'd7: my_line = line_7[frame_i];
            4'd8: my_line = line_8[frame_i];
            4'd9: my_line = line_9[frame_i];
            4'd10: my_line = line_10[frame_i];
            4'd11: my_line = line_11[frame_i];
            default: my_line = 'x;
        endcase
    end
    
    // Threshold must be shifted
    always_comb begin
        case (line_i)
            4'd0: my_thresh = threshold_9[frame_i];
            4'd1: my_thresh = threshold_10[frame_i];
            4'd2: my_thresh = threshold_11[frame_i];
            4'd3: my_thresh = threshold_0[frame_i];
            4'd4: my_thresh = threshold_1[frame_i];
            4'd5: my_thresh = threshold_2[frame_i];
            4'd6: my_thresh = threshold_3[frame_i];
            4'd7: my_thresh = threshold_4[frame_i];
            4'd8: my_thresh = threshold_5[frame_i];
            4'd9: my_thresh = threshold_6[frame_i];
            4'd10: my_thresh = threshold_7[frame_i];
            4'd11: my_thresh = threshold_8[frame_i];
            default: my_thresh = 'x;
        endcase
    end
    
logic [4*types::LINE_BITS-1:0] line_0 [32];
logic [types::THRESH_BITS-1:0] threshold_0 [32];
assign line_0[0] = {7'd22, 7'd17, 7'd80, 7'd17};
assign threshold_0[0] = 8'd58;
assign line_0[1] = {7'd19, 7'd15, 7'd76, 7'd19};
assign threshold_0[1] = 8'd57;
assign line_0[2] = {7'd17, 7'd14, 7'd70, 7'd21};
assign threshold_0[2] = 8'd53;
assign line_0[3] = {7'd17, 7'd12, 7'd63, 7'd22};
assign threshold_0[3] = 8'd47;
assign line_0[4] = {7'd18, 7'd10, 7'd56, 7'd21};
assign threshold_0[4] = 8'd40;
assign line_0[5] = {7'd20, 7'd9, 7'd49, 7'd20};
assign threshold_0[5] = 8'd31;
assign line_0[6] = {7'd24, 7'd8, 7'd43, 7'd17};
assign threshold_0[6] = 8'd21;
assign line_0[7] = {7'd29, 7'd8, 7'd38, 7'd14};
assign threshold_0[7] = 8'd11;
assign line_0[8] = {7'd35, 7'd10, 7'd35, 7'd10};
assign threshold_0[8] = 8'd0;
assign line_0[9] = {7'd34, 7'd7, 7'd41, 7'd13};
assign threshold_0[9] = 8'd9;
assign line_0[10] = {7'd34, 7'd4, 7'd46, 7'd18};
assign threshold_0[10] = 8'd18;
assign line_0[11] = {7'd36, 7'd3, 7'd51, 7'd23};
assign threshold_0[11] = 8'd25;
assign line_0[12] = {7'd39, 7'd3, 7'd55, 7'd30};
assign threshold_0[12] = 8'd31;
assign line_0[13] = {7'd43, 7'd4, 7'd57, 7'd37};
assign threshold_0[13] = 8'd36;
assign line_0[14] = {7'd46, 7'd7, 7'd57, 7'd45};
assign threshold_0[14] = 8'd40;
assign line_0[15] = {7'd49, 7'd11, 7'd55, 7'd52};
assign threshold_0[15] = 8'd41;
assign line_0[16] = {7'd51, 7'd17, 7'd50, 7'd59};
assign threshold_0[16] = 8'd42;
assign line_0[17] = {7'd51, 7'd23, 7'd45, 7'd64};
assign threshold_0[17] = 8'd41;
assign line_0[18] = {7'd49, 7'd29, 7'd38, 7'd67};
assign threshold_0[18] = 8'd40;
assign line_0[19] = {7'd45, 7'd35, 7'd31, 7'd69};
assign threshold_0[19] = 8'd37;
assign line_0[20] = {7'd40, 7'd41, 7'd24, 7'd68};
assign threshold_0[20] = 8'd31;
assign line_0[21] = {7'd34, 7'd45, 7'd19, 7'd66};
assign threshold_0[21] = 8'd26;
assign line_0[22] = {7'd27, 7'd48, 7'd14, 7'd61};
assign threshold_0[22] = 8'd18;
assign line_0[23] = {7'd19, 7'd49, 7'd12, 7'd56};
assign threshold_0[23] = 8'd10;
assign line_0[24] = {7'd13, 7'd49, 7'd13, 7'd49};
assign threshold_0[24] = 8'd0;
assign line_0[25] = {7'd16, 7'd42, 7'd7, 7'd47};
assign threshold_0[25] = 8'd10;
assign line_0[26] = {7'd21, 7'd35, 7'd3, 7'd44};
assign threshold_0[26] = 8'd20;
assign line_0[27] = {7'd29, 7'd29, 7'd1, 7'd40};
assign threshold_0[27] = 8'd30;
assign line_0[28] = {7'd38, 7'd23, 7'd1, 7'd35};
assign threshold_0[28] = 8'd39;
assign line_0[29] = {7'd49, 7'd19, 7'd3, 7'd29};
assign threshold_0[29] = 8'd47;
assign line_0[30] = {7'd60, 7'd17, 7'd7, 7'd25};
assign threshold_0[30] = 8'd54;
assign line_0[31] = {7'd70, 7'd16, 7'd14, 7'd20};
assign threshold_0[31] = 8'd56;
logic [4*types::LINE_BITS-1:0] line_1 [32];
logic [types::THRESH_BITS-1:0] threshold_1 [32];
assign line_1[0] = {7'd80, 7'd17, 7'd80, 7'd17};
assign threshold_1[0] = 8'd0;
assign line_1[1] = {7'd87, 7'd18, 7'd76, 7'd19};
assign threshold_1[1] = 8'd11;
assign line_1[2] = {7'd93, 7'd20, 7'd70, 7'd21};
assign threshold_1[2] = 8'd23;
assign line_1[3] = {7'd63, 7'd22, 7'd96, 7'd23};
assign threshold_1[3] = 8'd33;
assign line_1[4] = {7'd56, 7'd21, 7'd97, 7'd25};
assign threshold_1[4] = 8'd41;
assign line_1[5] = {7'd49, 7'd20, 7'd97, 7'd27};
assign threshold_1[5] = 8'd49;
assign line_1[6] = {7'd43, 7'd17, 7'd95, 7'd27};
assign threshold_1[6] = 8'd53;
assign line_1[7] = {7'd38, 7'd14, 7'd92, 7'd27};
assign threshold_1[7] = 8'd56;
assign line_1[8] = {7'd35, 7'd10, 7'd88, 7'd26};
assign threshold_1[8] = 8'd55;
assign line_1[9] = {7'd34, 7'd7, 7'd85, 7'd24};
assign threshold_1[9] = 8'd54;
assign line_1[10] = {7'd34, 7'd4, 7'd83, 7'd22};
assign threshold_1[10] = 8'd52;
assign line_1[11] = {7'd36, 7'd3, 7'd82, 7'd19};
assign threshold_1[11] = 8'd49;
assign line_1[12] = {7'd39, 7'd3, 7'd82, 7'd16};
assign threshold_1[12] = 8'd45;
assign line_1[13] = {7'd43, 7'd4, 7'd83, 7'd15};
assign threshold_1[13] = 8'd41;
assign line_1[14] = {7'd46, 7'd7, 7'd86, 7'd14};
assign threshold_1[14] = 8'd41;
assign line_1[15] = {7'd49, 7'd11, 7'd89, 7'd14};
assign threshold_1[15] = 8'd40;
assign line_1[16] = {7'd51, 7'd17, 7'd92, 7'd17};
assign threshold_1[16] = 8'd41;
assign line_1[17] = {7'd94, 7'd20, 7'd51, 7'd23};
assign threshold_1[17] = 8'd43;
assign line_1[18] = {7'd95, 7'd25, 7'd49, 7'd29};
assign threshold_1[18] = 8'd46;
assign line_1[19] = {7'd95, 7'd32, 7'd45, 7'd35};
assign threshold_1[19] = 8'd50;
assign line_1[20] = {7'd93, 7'd39, 7'd40, 7'd41};
assign threshold_1[20] = 8'd53;
assign line_1[21] = {7'd34, 7'd45, 7'd89, 7'd46};
assign threshold_1[21] = 8'd55;
assign line_1[22] = {7'd27, 7'd48, 7'd83, 7'd53};
assign threshold_1[22] = 8'd56;
assign line_1[23] = {7'd19, 7'd49, 7'd75, 7'd60};
assign threshold_1[23] = 8'd57;
assign line_1[24] = {7'd13, 7'd49, 7'd66, 7'd65};
assign threshold_1[24] = 8'd55;
assign line_1[25] = {7'd7, 7'd47, 7'd56, 7'd69};
assign threshold_1[25] = 8'd54;
assign line_1[26] = {7'd3, 7'd44, 7'd47, 7'd71};
assign threshold_1[26] = 8'd52;
assign line_1[27] = {7'd1, 7'd40, 7'd37, 7'd71};
assign threshold_1[27] = 8'd48;
assign line_1[28] = {7'd1, 7'd35, 7'd30, 7'd70};
assign threshold_1[28] = 8'd45;
assign line_1[29] = {7'd3, 7'd29, 7'd24, 7'd68};
assign threshold_1[29] = 8'd44;
assign line_1[30] = {7'd7, 7'd25, 7'd21, 7'd65};
assign threshold_1[30] = 8'd42;
assign line_1[31] = {7'd14, 7'd20, 7'd20, 7'd62};
assign threshold_1[31] = 8'd42;
logic [4*types::LINE_BITS-1:0] line_2 [32];
logic [types::THRESH_BITS-1:0] threshold_2 [32];
assign line_2[0] = {7'd80, 7'd17, 7'd22, 7'd17};
assign threshold_2[0] = 8'd58;
assign line_2[1] = {7'd31, 7'd14, 7'd87, 7'd18};
assign threshold_2[1] = 8'd56;
assign line_2[2] = {7'd40, 7'd13, 7'd93, 7'd20};
assign threshold_2[2] = 8'd53;
assign line_2[3] = {7'd50, 7'd12, 7'd96, 7'd23};
assign threshold_2[3] = 8'd47;
assign line_2[4] = {7'd59, 7'd13, 7'd97, 7'd25};
assign threshold_2[4] = 8'd40;
assign line_2[5] = {7'd68, 7'd16, 7'd97, 7'd27};
assign threshold_2[5] = 8'd31;
assign line_2[6] = {7'd76, 7'd18, 7'd95, 7'd27};
assign threshold_2[6] = 8'd21;
assign line_2[7] = {7'd83, 7'd22, 7'd92, 7'd27};
assign threshold_2[7] = 8'd10;
assign line_2[8] = {7'd88, 7'd26, 7'd88, 7'd26};
assign threshold_2[8] = 8'd0;
assign line_2[9] = {7'd85, 7'd24, 7'd93, 7'd31};
assign threshold_2[9] = 8'd11;
assign line_2[10] = {7'd83, 7'd22, 7'd95, 7'd35};
assign threshold_2[10] = 8'd18;
assign line_2[11] = {7'd82, 7'd19, 7'd97, 7'd40};
assign threshold_2[11] = 8'd26;
assign line_2[12] = {7'd82, 7'd16, 7'd98, 7'd44};
assign threshold_2[12] = 8'd32;
assign line_2[13] = {7'd83, 7'd15, 7'd97, 7'd48};
assign threshold_2[13] = 8'd36;
assign line_2[14] = {7'd86, 7'd14, 7'd96, 7'd52};
assign threshold_2[14] = 8'd39;
assign line_2[15] = {7'd89, 7'd14, 7'd94, 7'd55};
assign threshold_2[15] = 8'd41;
assign line_2[16] = {7'd92, 7'd17, 7'd92, 7'd59};
assign threshold_2[16] = 8'd42;
assign line_2[17] = {7'd94, 7'd20, 7'd88, 7'd61};
assign threshold_2[17] = 8'd41;
assign line_2[18] = {7'd95, 7'd25, 7'd85, 7'd63};
assign threshold_2[18] = 8'd39;
assign line_2[19] = {7'd95, 7'd32, 7'd81, 7'd65};
assign threshold_2[19] = 8'd36;
assign line_2[20] = {7'd93, 7'd39, 7'd78, 7'd66};
assign threshold_2[20] = 8'd31;
assign line_2[21] = {7'd89, 7'd46, 7'd74, 7'd67};
assign threshold_2[21] = 8'd26;
assign line_2[22] = {7'd83, 7'd53, 7'd71, 7'd67};
assign threshold_2[22] = 8'd18;
assign line_2[23] = {7'd75, 7'd60, 7'd68, 7'd66};
assign threshold_2[23] = 8'd9;
assign line_2[24] = {7'd66, 7'd65, 7'd66, 7'd65};
assign threshold_2[24] = 8'd0;
assign line_2[25] = {7'd65, 7'd64, 7'd56, 7'd69};
assign threshold_2[25] = 8'd10;
assign line_2[26] = {7'd65, 7'd62, 7'd47, 7'd71};
assign threshold_2[26] = 8'd20;
assign line_2[27] = {7'd66, 7'd60, 7'd37, 7'd71};
assign threshold_2[27] = 8'd31;
assign line_2[28] = {7'd68, 7'd59, 7'd30, 7'd70};
assign threshold_2[28] = 8'd40;
assign line_2[29] = {7'd70, 7'd58, 7'd24, 7'd68};
assign threshold_2[29] = 8'd47;
assign line_2[30] = {7'd73, 7'd58, 7'd21, 7'd65};
assign threshold_2[30] = 8'd52;
assign line_2[31] = {7'd76, 7'd58, 7'd20, 7'd62};
assign threshold_2[31] = 8'd56;
logic [4*types::LINE_BITS-1:0] line_3 [32];
logic [types::THRESH_BITS-1:0] threshold_3 [32];
assign line_3[0] = {7'd22, 7'd17, 7'd22, 7'd17};
assign threshold_3[0] = 8'd0;
assign line_3[1] = {7'd31, 7'd14, 7'd19, 7'd15};
assign threshold_3[1] = 8'd12;
assign line_3[2] = {7'd40, 7'd13, 7'd17, 7'd14};
assign threshold_3[2] = 8'd23;
assign line_3[3] = {7'd50, 7'd12, 7'd17, 7'd12};
assign threshold_3[3] = 8'd33;
assign line_3[4] = {7'd18, 7'd10, 7'd59, 7'd13};
assign threshold_3[4] = 8'd41;
assign line_3[5] = {7'd20, 7'd9, 7'd68, 7'd16};
assign threshold_3[5] = 8'd49;
assign line_3[6] = {7'd24, 7'd8, 7'd76, 7'd18};
assign threshold_3[6] = 8'd53;
assign line_3[7] = {7'd29, 7'd8, 7'd83, 7'd22};
assign threshold_3[7] = 8'd56;
assign line_3[8] = {7'd35, 7'd10, 7'd88, 7'd26};
assign threshold_3[8] = 8'd55;
assign line_3[9] = {7'd41, 7'd13, 7'd93, 7'd31};
assign threshold_3[9] = 8'd55;
assign line_3[10] = {7'd46, 7'd18, 7'd95, 7'd35};
assign threshold_3[10] = 8'd52;
assign line_3[11] = {7'd51, 7'd23, 7'd97, 7'd40};
assign threshold_3[11] = 8'd49;
assign line_3[12] = {7'd55, 7'd30, 7'd98, 7'd44};
assign threshold_3[12] = 8'd45;
assign line_3[13] = {7'd57, 7'd37, 7'd97, 7'd48};
assign threshold_3[13] = 8'd41;
assign line_3[14] = {7'd57, 7'd45, 7'd96, 7'd52};
assign threshold_3[14] = 8'd40;
assign line_3[15] = {7'd55, 7'd52, 7'd94, 7'd55};
assign threshold_3[15] = 8'd39;
assign line_3[16] = {7'd92, 7'd59, 7'd50, 7'd59};
assign threshold_3[16] = 8'd42;
assign line_3[17] = {7'd88, 7'd61, 7'd45, 7'd64};
assign threshold_3[17] = 8'd43;
assign line_3[18] = {7'd85, 7'd63, 7'd38, 7'd67};
assign threshold_3[18] = 8'd47;
assign line_3[19] = {7'd81, 7'd65, 7'd31, 7'd69};
assign threshold_3[19] = 8'd50;
assign line_3[20] = {7'd78, 7'd66, 7'd24, 7'd68};
assign threshold_3[20] = 8'd54;
assign line_3[21] = {7'd19, 7'd66, 7'd74, 7'd67};
assign threshold_3[21] = 8'd55;
assign line_3[22] = {7'd14, 7'd61, 7'd71, 7'd67};
assign threshold_3[22] = 8'd57;
assign line_3[23] = {7'd12, 7'd56, 7'd68, 7'd66};
assign threshold_3[23] = 8'd57;
assign line_3[24] = {7'd13, 7'd49, 7'd66, 7'd65};
assign threshold_3[24] = 8'd55;
assign line_3[25] = {7'd16, 7'd42, 7'd65, 7'd64};
assign threshold_3[25] = 8'd54;
assign line_3[26] = {7'd21, 7'd35, 7'd65, 7'd62};
assign threshold_3[26] = 8'd52;
assign line_3[27] = {7'd29, 7'd29, 7'd66, 7'd60};
assign threshold_3[27] = 8'd48;
assign line_3[28] = {7'd38, 7'd23, 7'd68, 7'd59};
assign threshold_3[28] = 8'd47;
assign line_3[29] = {7'd49, 7'd19, 7'd70, 7'd58};
assign threshold_3[29] = 8'd44;
assign line_3[30] = {7'd60, 7'd17, 7'd73, 7'd58};
assign threshold_3[30] = 8'd43;
assign line_3[31] = {7'd70, 7'd16, 7'd76, 7'd58};
assign threshold_3[31] = 8'd42;
logic [4*types::LINE_BITS-1:0] line_4 [32];
logic [types::THRESH_BITS-1:0] threshold_4 [32];
assign line_4[0] = {7'd22, 7'd17, 7'd22, 7'd59};
assign threshold_4[0] = 8'd42;
assign line_4[1] = {7'd19, 7'd15, 7'd14, 7'd57};
assign threshold_4[1] = 8'd42;
assign line_4[2] = {7'd17, 7'd14, 7'd8, 7'd55};
assign threshold_4[2] = 8'd42;
assign line_4[3] = {7'd17, 7'd12, 7'd5, 7'd52};
assign threshold_4[3] = 8'd42;
assign line_4[4] = {7'd18, 7'd10, 7'd4, 7'd50};
assign threshold_4[4] = 8'd42;
assign line_4[5] = {7'd20, 7'd9, 7'd4, 7'd48};
assign threshold_4[5] = 8'd42;
assign line_4[6] = {7'd24, 7'd8, 7'd6, 7'd48};
assign threshold_4[6] = 8'd44;
assign line_4[7] = {7'd29, 7'd8, 7'd9, 7'd48};
assign threshold_4[7] = 8'd45;
assign line_4[8] = {7'd35, 7'd10, 7'd13, 7'd49};
assign threshold_4[8] = 8'd45;
assign line_4[9] = {7'd41, 7'd13, 7'd16, 7'd51};
assign threshold_4[9] = 8'd45;
assign line_4[10] = {7'd46, 7'd18, 7'd18, 7'd53};
assign threshold_4[10] = 8'd45;
assign line_4[11] = {7'd51, 7'd23, 7'd19, 7'd56};
assign threshold_4[11] = 8'd46;
assign line_4[12] = {7'd55, 7'd30, 7'd19, 7'd59};
assign threshold_4[12] = 8'd46;
assign line_4[13] = {7'd57, 7'd37, 7'd18, 7'd60};
assign threshold_4[13] = 8'd45;
assign line_4[14] = {7'd57, 7'd45, 7'd15, 7'd61};
assign threshold_4[14] = 8'd45;
assign line_4[15] = {7'd55, 7'd52, 7'd12, 7'd61};
assign threshold_4[15] = 8'd44;
assign line_4[16] = {7'd9, 7'd58, 7'd50, 7'd59};
assign threshold_4[16] = 8'd41;
assign line_4[17] = {7'd7, 7'd55, 7'd45, 7'd64};
assign threshold_4[17] = 8'd39;
assign line_4[18] = {7'd6, 7'd50, 7'd38, 7'd67};
assign threshold_4[18] = 8'd36;
assign line_4[19] = {7'd6, 7'd43, 7'd31, 7'd69};
assign threshold_4[19] = 8'd36;
assign line_4[20] = {7'd8, 7'd36, 7'd24, 7'd68};
assign threshold_4[20] = 8'd36;
assign line_4[21] = {7'd12, 7'd29, 7'd19, 7'd66};
assign threshold_4[21] = 8'd38;
assign line_4[22] = {7'd18, 7'd22, 7'd14, 7'd61};
assign threshold_4[22] = 8'd39;
assign line_4[23] = {7'd26, 7'd15, 7'd12, 7'd56};
assign threshold_4[23] = 8'd43;
assign line_4[24] = {7'd35, 7'd10, 7'd13, 7'd49};
assign threshold_4[24] = 8'd45;
assign line_4[25] = {7'd45, 7'd6, 7'd16, 7'd42};
assign threshold_4[25] = 8'd46;
assign line_4[26] = {7'd54, 7'd4, 7'd21, 7'd35};
assign threshold_4[26] = 8'd45;
assign line_4[27] = {7'd64, 7'd4, 7'd29, 7'd29};
assign threshold_4[27] = 8'd43;
assign line_4[28] = {7'd71, 7'd5, 7'd38, 7'd23};
assign threshold_4[28] = 8'd38;
assign line_4[29] = {7'd77, 7'd7, 7'd49, 7'd19};
assign threshold_4[29] = 8'd30;
assign line_4[30] = {7'd80, 7'd10, 7'd60, 7'd17};
assign threshold_4[30] = 8'd21;
assign line_4[31] = {7'd81, 7'd13, 7'd70, 7'd16};
assign threshold_4[31] = 8'd11;
logic [4*types::LINE_BITS-1:0] line_5 [32];
logic [types::THRESH_BITS-1:0] threshold_5 [32];
assign line_5[0] = {7'd80, 7'd17, 7'd80, 7'd59};
assign threshold_5[0] = 8'd42;
assign line_5[1] = {7'd76, 7'd19, 7'd70, 7'd61};
assign threshold_5[1] = 8'd42;
assign line_5[2] = {7'd70, 7'd21, 7'd61, 7'd62};
assign threshold_5[2] = 8'd42;
assign line_5[3] = {7'd63, 7'd22, 7'd51, 7'd63};
assign threshold_5[3] = 8'd43;
assign line_5[4] = {7'd56, 7'd21, 7'd42, 7'd62};
assign threshold_5[4] = 8'd43;
assign line_5[5] = {7'd49, 7'd20, 7'd33, 7'd59};
assign threshold_5[5] = 8'd42;
assign line_5[6] = {7'd43, 7'd17, 7'd25, 7'd57};
assign threshold_5[6] = 8'd44;
assign line_5[7] = {7'd38, 7'd14, 7'd18, 7'd53};
assign threshold_5[7] = 8'd44;
assign line_5[8] = {7'd35, 7'd10, 7'd13, 7'd49};
assign threshold_5[8] = 8'd45;
assign line_5[9] = {7'd34, 7'd7, 7'd8, 7'd44};
assign threshold_5[9] = 8'd45;
assign line_5[10] = {7'd34, 7'd4, 7'd6, 7'd40};
assign threshold_5[10] = 8'd46;
assign line_5[11] = {7'd36, 7'd3, 7'd4, 7'd35};
assign threshold_5[11] = 8'd45;
assign line_5[12] = {7'd39, 7'd3, 7'd3, 7'd31};
assign threshold_5[12] = 8'd46;
assign line_5[13] = {7'd43, 7'd4, 7'd4, 7'd27};
assign threshold_5[13] = 8'd45;
assign line_5[14] = {7'd46, 7'd7, 7'd5, 7'd23};
assign threshold_5[14] = 8'd44;
assign line_5[15] = {7'd49, 7'd11, 7'd7, 7'd20};
assign threshold_5[15] = 8'd43;
assign line_5[16] = {7'd9, 7'd16, 7'd51, 7'd17};
assign threshold_5[16] = 8'd42;
assign line_5[17] = {7'd13, 7'd14, 7'd51, 7'd23};
assign threshold_5[17] = 8'd39;
assign line_5[18] = {7'd16, 7'd12, 7'd49, 7'd29};
assign threshold_5[18] = 8'd37;
assign line_5[19] = {7'd20, 7'd10, 7'd45, 7'd35};
assign threshold_5[19] = 8'd35;
assign line_5[20] = {7'd23, 7'd9, 7'd40, 7'd41};
assign threshold_5[20] = 8'd36;
assign line_5[21] = {7'd27, 7'd8, 7'd34, 7'd45};
assign threshold_5[21] = 8'd38;
assign line_5[22] = {7'd30, 7'd8, 7'd27, 7'd48};
assign threshold_5[22] = 8'd40;
assign line_5[23] = {7'd33, 7'd9, 7'd19, 7'd49};
assign threshold_5[23] = 8'd42;
assign line_5[24] = {7'd35, 7'd10, 7'd13, 7'd49};
assign threshold_5[24] = 8'd45;
assign line_5[25] = {7'd36, 7'd11, 7'd7, 7'd47};
assign threshold_5[25] = 8'd46;
assign line_5[26] = {7'd36, 7'd13, 7'd3, 7'd44};
assign threshold_5[26] = 8'd45;
assign line_5[27] = {7'd35, 7'd15, 7'd1, 7'd40};
assign threshold_5[27] = 8'd42;
assign line_5[28] = {7'd33, 7'd16, 7'd1, 7'd35};
assign threshold_5[28] = 8'd37;
assign line_5[29] = {7'd31, 7'd17, 7'd3, 7'd29};
assign threshold_5[29] = 8'd30;
assign line_5[30] = {7'd28, 7'd17, 7'd7, 7'd25};
assign threshold_5[30] = 8'd22;
assign line_5[31] = {7'd25, 7'd17, 7'd14, 7'd20};
assign threshold_5[31] = 8'd11;
logic [4*types::LINE_BITS-1:0] line_6 [32];
logic [types::THRESH_BITS-1:0] threshold_6 [32];
assign line_6[0] = {7'd22, 7'd17, 7'd22, 7'd59};
assign threshold_6[0] = 8'd42;
assign line_6[1] = {7'd31, 7'd14, 7'd25, 7'd56};
assign threshold_6[1] = 8'd42;
assign line_6[2] = {7'd40, 7'd13, 7'd31, 7'd54};
assign threshold_6[2] = 8'd42;
assign line_6[3] = {7'd50, 7'd12, 7'd38, 7'd53};
assign threshold_6[3] = 8'd43;
assign line_6[4] = {7'd59, 7'd13, 7'd45, 7'd54};
assign threshold_6[4] = 8'd43;
assign line_6[5] = {7'd68, 7'd16, 7'd52, 7'd55};
assign threshold_6[5] = 8'd42;
assign line_6[6] = {7'd76, 7'd18, 7'd58, 7'd58};
assign threshold_6[6] = 8'd44;
assign line_6[7] = {7'd83, 7'd22, 7'd63, 7'd61};
assign threshold_6[7] = 8'd44;
assign line_6[8] = {7'd88, 7'd26, 7'd66, 7'd65};
assign threshold_6[8] = 8'd45;
assign line_6[9] = {7'd93, 7'd31, 7'd67, 7'd68};
assign threshold_6[9] = 8'd45;
assign line_6[10] = {7'd95, 7'd35, 7'd67, 7'd71};
assign threshold_6[10] = 8'd46;
assign line_6[11] = {7'd97, 7'd40, 7'd65, 7'd72};
assign threshold_6[11] = 8'd45;
assign line_6[12] = {7'd98, 7'd44, 7'd62, 7'd72};
assign threshold_6[12] = 8'd46;
assign line_6[13] = {7'd97, 7'd48, 7'd58, 7'd71};
assign threshold_6[13] = 8'd45;
assign line_6[14] = {7'd96, 7'd52, 7'd55, 7'd68};
assign threshold_6[14] = 8'd44;
assign line_6[15] = {7'd94, 7'd55, 7'd52, 7'd64};
assign threshold_6[15] = 8'd43;
assign line_6[16] = {7'd51, 7'd58, 7'd92, 7'd59};
assign threshold_6[16] = 8'd41;
assign line_6[17] = {7'd50, 7'd52, 7'd88, 7'd61};
assign threshold_6[17] = 8'd39;
assign line_6[18] = {7'd52, 7'd46, 7'd85, 7'd63};
assign threshold_6[18] = 8'd37;
assign line_6[19] = {7'd56, 7'd40, 7'd81, 7'd65};
assign threshold_6[19] = 8'd35;
assign line_6[20] = {7'd61, 7'd34, 7'd78, 7'd66};
assign threshold_6[20] = 8'd36;
assign line_6[21] = {7'd67, 7'd30, 7'd74, 7'd67};
assign threshold_6[21] = 8'd38;
assign line_6[22] = {7'd74, 7'd27, 7'd71, 7'd67};
assign threshold_6[22] = 8'd40;
assign line_6[23] = {7'd82, 7'd26, 7'd68, 7'd66};
assign threshold_6[23] = 8'd42;
assign line_6[24] = {7'd88, 7'd26, 7'd66, 7'd65};
assign threshold_6[24] = 8'd45;
assign line_6[25] = {7'd94, 7'd28, 7'd65, 7'd64};
assign threshold_6[25] = 8'd46;
assign line_6[26] = {7'd98, 7'd31, 7'd65, 7'd62};
assign threshold_6[26] = 8'd45;
assign line_6[27] = {7'd100, 7'd35, 7'd66, 7'd60};
assign threshold_6[27] = 8'd42;
assign line_6[28] = {7'd100, 7'd40, 7'd68, 7'd59};
assign threshold_6[28] = 8'd37;
assign line_6[29] = {7'd98, 7'd46, 7'd70, 7'd58};
assign threshold_6[29] = 8'd30;
assign line_6[30] = {7'd94, 7'd50, 7'd73, 7'd58};
assign threshold_6[30] = 8'd22;
assign line_6[31] = {7'd87, 7'd55, 7'd76, 7'd58};
assign threshold_6[31] = 8'd11;
logic [4*types::LINE_BITS-1:0] line_7 [32];
logic [types::THRESH_BITS-1:0] threshold_7 [32];
assign line_7[0] = {7'd80, 7'd17, 7'd80, 7'd59};
assign threshold_7[0] = 8'd42;
assign line_7[1] = {7'd87, 7'd18, 7'd82, 7'd60};
assign threshold_7[1] = 8'd42;
assign line_7[2] = {7'd93, 7'd20, 7'd84, 7'd61};
assign threshold_7[2] = 8'd42;
assign line_7[3] = {7'd96, 7'd23, 7'd84, 7'd63};
assign threshold_7[3] = 8'd42;
assign line_7[4] = {7'd97, 7'd25, 7'd83, 7'd65};
assign threshold_7[4] = 8'd42;
assign line_7[5] = {7'd97, 7'd27, 7'd81, 7'd66};
assign threshold_7[5] = 8'd42;
assign line_7[6] = {7'd95, 7'd27, 7'd77, 7'd67};
assign threshold_7[6] = 8'd44;
assign line_7[7] = {7'd92, 7'd27, 7'd72, 7'd67};
assign threshold_7[7] = 8'd45;
assign line_7[8] = {7'd88, 7'd26, 7'd66, 7'd65};
assign threshold_7[8] = 8'd45;
assign line_7[9] = {7'd85, 7'd24, 7'd60, 7'd62};
assign threshold_7[9] = 8'd45;
assign line_7[10] = {7'd83, 7'd22, 7'd55, 7'd57};
assign threshold_7[10] = 8'd45;
assign line_7[11] = {7'd82, 7'd19, 7'd50, 7'd52};
assign threshold_7[11] = 8'd46;
assign line_7[12] = {7'd82, 7'd16, 7'd46, 7'd45};
assign threshold_7[12] = 8'd46;
assign line_7[13] = {7'd83, 7'd15, 7'd44, 7'd38};
assign threshold_7[13] = 8'd45;
assign line_7[14] = {7'd86, 7'd14, 7'd44, 7'd30};
assign threshold_7[14] = 8'd45;
assign line_7[15] = {7'd89, 7'd14, 7'd46, 7'd23};
assign threshold_7[15] = 8'd44;
assign line_7[16] = {7'd51, 7'd16, 7'd92, 7'd17};
assign threshold_7[16] = 8'd41;
assign line_7[17] = {7'd56, 7'd11, 7'd94, 7'd20};
assign threshold_7[17] = 8'd39;
assign line_7[18] = {7'd63, 7'd8, 7'd95, 7'd25};
assign threshold_7[18] = 8'd36;
assign line_7[19] = {7'd70, 7'd6, 7'd95, 7'd32};
assign threshold_7[19] = 8'd36;
assign line_7[20] = {7'd77, 7'd7, 7'd93, 7'd39};
assign threshold_7[20] = 8'd36;
assign line_7[21] = {7'd82, 7'd9, 7'd89, 7'd46};
assign threshold_7[21] = 8'd38;
assign line_7[22] = {7'd87, 7'd14, 7'd83, 7'd53};
assign threshold_7[22] = 8'd39;
assign line_7[23] = {7'd89, 7'd19, 7'd75, 7'd60};
assign threshold_7[23] = 8'd43;
assign line_7[24] = {7'd88, 7'd26, 7'd66, 7'd65};
assign threshold_7[24] = 8'd45;
assign line_7[25] = {7'd85, 7'd33, 7'd56, 7'd69};
assign threshold_7[25] = 8'd46;
assign line_7[26] = {7'd80, 7'd40, 7'd47, 7'd71};
assign threshold_7[26] = 8'd45;
assign line_7[27] = {7'd72, 7'd46, 7'd37, 7'd71};
assign threshold_7[27] = 8'd43;
assign line_7[28] = {7'd63, 7'd52, 7'd30, 7'd70};
assign threshold_7[28] = 8'd38;
assign line_7[29] = {7'd52, 7'd56, 7'd24, 7'd68};
assign threshold_7[29] = 8'd30;
assign line_7[30] = {7'd41, 7'd58, 7'd21, 7'd65};
assign threshold_7[30] = 8'd21;
assign line_7[31] = {7'd31, 7'd59, 7'd20, 7'd62};
assign threshold_7[31] = 8'd11;
logic [4*types::LINE_BITS-1:0] line_8 [32];
logic [types::THRESH_BITS-1:0] threshold_8 [32];
assign line_8[0] = {7'd22, 7'd59, 7'd80, 7'd59};
assign threshold_8[0] = 8'd58;
assign line_8[1] = {7'd14, 7'd57, 7'd70, 7'd61};
assign threshold_8[1] = 8'd56;
assign line_8[2] = {7'd8, 7'd55, 7'd61, 7'd62};
assign threshold_8[2] = 8'd53;
assign line_8[3] = {7'd5, 7'd52, 7'd51, 7'd63};
assign threshold_8[3] = 8'd47;
assign line_8[4] = {7'd4, 7'd50, 7'd42, 7'd62};
assign threshold_8[4] = 8'd40;
assign line_8[5] = {7'd4, 7'd48, 7'd33, 7'd59};
assign threshold_8[5] = 8'd31;
assign line_8[6] = {7'd6, 7'd48, 7'd25, 7'd57};
assign threshold_8[6] = 8'd21;
assign line_8[7] = {7'd9, 7'd48, 7'd18, 7'd53};
assign threshold_8[7] = 8'd10;
assign line_8[8] = {7'd13, 7'd49, 7'd13, 7'd49};
assign threshold_8[8] = 8'd0;
assign line_8[9] = {7'd8, 7'd44, 7'd16, 7'd51};
assign threshold_8[9] = 8'd11;
assign line_8[10] = {7'd6, 7'd40, 7'd18, 7'd53};
assign threshold_8[10] = 8'd18;
assign line_8[11] = {7'd4, 7'd35, 7'd19, 7'd56};
assign threshold_8[11] = 8'd26;
assign line_8[12] = {7'd3, 7'd31, 7'd19, 7'd59};
assign threshold_8[12] = 8'd32;
assign line_8[13] = {7'd4, 7'd27, 7'd18, 7'd60};
assign threshold_8[13] = 8'd36;
assign line_8[14] = {7'd5, 7'd23, 7'd15, 7'd61};
assign threshold_8[14] = 8'd39;
assign line_8[15] = {7'd7, 7'd20, 7'd12, 7'd61};
assign threshold_8[15] = 8'd41;
assign line_8[16] = {7'd9, 7'd16, 7'd9, 7'd58};
assign threshold_8[16] = 8'd42;
assign line_8[17] = {7'd13, 7'd14, 7'd7, 7'd55};
assign threshold_8[17] = 8'd41;
assign line_8[18] = {7'd16, 7'd12, 7'd6, 7'd50};
assign threshold_8[18] = 8'd39;
assign line_8[19] = {7'd20, 7'd10, 7'd6, 7'd43};
assign threshold_8[19] = 8'd36;
assign line_8[20] = {7'd23, 7'd9, 7'd8, 7'd36};
assign threshold_8[20] = 8'd31;
assign line_8[21] = {7'd27, 7'd8, 7'd12, 7'd29};
assign threshold_8[21] = 8'd26;
assign line_8[22] = {7'd30, 7'd8, 7'd18, 7'd22};
assign threshold_8[22] = 8'd18;
assign line_8[23] = {7'd33, 7'd9, 7'd26, 7'd15};
assign threshold_8[23] = 8'd9;
assign line_8[24] = {7'd35, 7'd10, 7'd35, 7'd10};
assign threshold_8[24] = 8'd0;
assign line_8[25] = {7'd45, 7'd6, 7'd36, 7'd11};
assign threshold_8[25] = 8'd10;
assign line_8[26] = {7'd54, 7'd4, 7'd36, 7'd13};
assign threshold_8[26] = 8'd20;
assign line_8[27] = {7'd64, 7'd4, 7'd35, 7'd15};
assign threshold_8[27] = 8'd31;
assign line_8[28] = {7'd71, 7'd5, 7'd33, 7'd16};
assign threshold_8[28] = 8'd40;
assign line_8[29] = {7'd77, 7'd7, 7'd31, 7'd17};
assign threshold_8[29] = 8'd47;
assign line_8[30] = {7'd80, 7'd10, 7'd28, 7'd17};
assign threshold_8[30] = 8'd52;
assign line_8[31] = {7'd81, 7'd13, 7'd25, 7'd17};
assign threshold_8[31] = 8'd56;
logic [4*types::LINE_BITS-1:0] line_9 [32];
logic [types::THRESH_BITS-1:0] threshold_9 [32];
assign line_9[0] = {7'd80, 7'd59, 7'd80, 7'd59};
assign threshold_9[0] = 8'd0;
assign line_9[1] = {7'd82, 7'd60, 7'd70, 7'd61};
assign threshold_9[1] = 8'd12;
assign line_9[2] = {7'd84, 7'd61, 7'd61, 7'd62};
assign threshold_9[2] = 8'd23;
assign line_9[3] = {7'd51, 7'd63, 7'd84, 7'd63};
assign threshold_9[3] = 8'd33;
assign line_9[4] = {7'd42, 7'd62, 7'd83, 7'd65};
assign threshold_9[4] = 8'd41;
assign line_9[5] = {7'd33, 7'd59, 7'd81, 7'd66};
assign threshold_9[5] = 8'd49;
assign line_9[6] = {7'd25, 7'd57, 7'd77, 7'd67};
assign threshold_9[6] = 8'd53;
assign line_9[7] = {7'd18, 7'd53, 7'd72, 7'd67};
assign threshold_9[7] = 8'd56;
assign line_9[8] = {7'd13, 7'd49, 7'd66, 7'd65};
assign threshold_9[8] = 8'd55;
assign line_9[9] = {7'd8, 7'd44, 7'd60, 7'd62};
assign threshold_9[9] = 8'd55;
assign line_9[10] = {7'd6, 7'd40, 7'd55, 7'd57};
assign threshold_9[10] = 8'd52;
assign line_9[11] = {7'd4, 7'd35, 7'd50, 7'd52};
assign threshold_9[11] = 8'd49;
assign line_9[12] = {7'd3, 7'd31, 7'd46, 7'd45};
assign threshold_9[12] = 8'd45;
assign line_9[13] = {7'd4, 7'd27, 7'd44, 7'd38};
assign threshold_9[13] = 8'd41;
assign line_9[14] = {7'd5, 7'd23, 7'd44, 7'd30};
assign threshold_9[14] = 8'd40;
assign line_9[15] = {7'd7, 7'd20, 7'd46, 7'd23};
assign threshold_9[15] = 8'd39;
assign line_9[16] = {7'd9, 7'd16, 7'd51, 7'd16};
assign threshold_9[16] = 8'd42;
assign line_9[17] = {7'd56, 7'd11, 7'd13, 7'd14};
assign threshold_9[17] = 8'd43;
assign line_9[18] = {7'd63, 7'd8, 7'd16, 7'd12};
assign threshold_9[18] = 8'd47;
assign line_9[19] = {7'd70, 7'd6, 7'd20, 7'd10};
assign threshold_9[19] = 8'd50;
assign line_9[20] = {7'd77, 7'd7, 7'd23, 7'd9};
assign threshold_9[20] = 8'd54;
assign line_9[21] = {7'd27, 7'd8, 7'd82, 7'd9};
assign threshold_9[21] = 8'd55;
assign line_9[22] = {7'd30, 7'd8, 7'd87, 7'd14};
assign threshold_9[22] = 8'd57;
assign line_9[23] = {7'd33, 7'd9, 7'd89, 7'd19};
assign threshold_9[23] = 8'd57;
assign line_9[24] = {7'd35, 7'd10, 7'd88, 7'd26};
assign threshold_9[24] = 8'd55;
assign line_9[25] = {7'd36, 7'd11, 7'd85, 7'd33};
assign threshold_9[25] = 8'd54;
assign line_9[26] = {7'd36, 7'd13, 7'd80, 7'd40};
assign threshold_9[26] = 8'd52;
assign line_9[27] = {7'd35, 7'd15, 7'd72, 7'd46};
assign threshold_9[27] = 8'd48;
assign line_9[28] = {7'd33, 7'd16, 7'd63, 7'd52};
assign threshold_9[28] = 8'd47;
assign line_9[29] = {7'd31, 7'd17, 7'd52, 7'd56};
assign threshold_9[29] = 8'd44;
assign line_9[30] = {7'd28, 7'd17, 7'd41, 7'd58};
assign threshold_9[30] = 8'd43;
assign line_9[31] = {7'd25, 7'd17, 7'd31, 7'd59};
assign threshold_9[31] = 8'd42;
logic [4*types::LINE_BITS-1:0] line_10 [32];
logic [types::THRESH_BITS-1:0] threshold_10 [32];
assign line_10[0] = {7'd80, 7'd59, 7'd22, 7'd59};
assign threshold_10[0] = 8'd58;
assign line_10[1] = {7'd25, 7'd56, 7'd82, 7'd60};
assign threshold_10[1] = 8'd57;
assign line_10[2] = {7'd31, 7'd54, 7'd84, 7'd61};
assign threshold_10[2] = 8'd53;
assign line_10[3] = {7'd38, 7'd53, 7'd84, 7'd63};
assign threshold_10[3] = 8'd47;
assign line_10[4] = {7'd45, 7'd54, 7'd83, 7'd65};
assign threshold_10[4] = 8'd40;
assign line_10[5] = {7'd52, 7'd55, 7'd81, 7'd66};
assign threshold_10[5] = 8'd31;
assign line_10[6] = {7'd58, 7'd58, 7'd77, 7'd67};
assign threshold_10[6] = 8'd21;
assign line_10[7] = {7'd63, 7'd61, 7'd72, 7'd67};
assign threshold_10[7] = 8'd11;
assign line_10[8] = {7'd66, 7'd65, 7'd66, 7'd65};
assign threshold_10[8] = 8'd0;
assign line_10[9] = {7'd60, 7'd62, 7'd67, 7'd68};
assign threshold_10[9] = 8'd9;
assign line_10[10] = {7'd55, 7'd57, 7'd67, 7'd71};
assign threshold_10[10] = 8'd18;
assign line_10[11] = {7'd50, 7'd52, 7'd65, 7'd72};
assign threshold_10[11] = 8'd25;
assign line_10[12] = {7'd46, 7'd45, 7'd62, 7'd72};
assign threshold_10[12] = 8'd31;
assign line_10[13] = {7'd44, 7'd38, 7'd58, 7'd71};
assign threshold_10[13] = 8'd36;
assign line_10[14] = {7'd44, 7'd30, 7'd55, 7'd68};
assign threshold_10[14] = 8'd40;
assign line_10[15] = {7'd46, 7'd23, 7'd52, 7'd64};
assign threshold_10[15] = 8'd41;
assign line_10[16] = {7'd51, 7'd16, 7'd51, 7'd58};
assign threshold_10[16] = 8'd42;
assign line_10[17] = {7'd56, 7'd11, 7'd50, 7'd52};
assign threshold_10[17] = 8'd41;
assign line_10[18] = {7'd63, 7'd8, 7'd52, 7'd46};
assign threshold_10[18] = 8'd40;
assign line_10[19] = {7'd70, 7'd6, 7'd56, 7'd40};
assign threshold_10[19] = 8'd37;
assign line_10[20] = {7'd77, 7'd7, 7'd61, 7'd34};
assign threshold_10[20] = 8'd31;
assign line_10[21] = {7'd82, 7'd9, 7'd67, 7'd30};
assign threshold_10[21] = 8'd26;
assign line_10[22] = {7'd87, 7'd14, 7'd74, 7'd27};
assign threshold_10[22] = 8'd18;
assign line_10[23] = {7'd89, 7'd19, 7'd82, 7'd26};
assign threshold_10[23] = 8'd10;
assign line_10[24] = {7'd88, 7'd26, 7'd88, 7'd26};
assign threshold_10[24] = 8'd0;
assign line_10[25] = {7'd94, 7'd28, 7'd85, 7'd33};
assign threshold_10[25] = 8'd10;
assign line_10[26] = {7'd98, 7'd31, 7'd80, 7'd40};
assign threshold_10[26] = 8'd20;
assign line_10[27] = {7'd100, 7'd35, 7'd72, 7'd46};
assign threshold_10[27] = 8'd30;
assign line_10[28] = {7'd100, 7'd40, 7'd63, 7'd52};
assign threshold_10[28] = 8'd39;
assign line_10[29] = {7'd98, 7'd46, 7'd52, 7'd56};
assign threshold_10[29] = 8'd47;
assign line_10[30] = {7'd94, 7'd50, 7'd41, 7'd58};
assign threshold_10[30] = 8'd54;
assign line_10[31] = {7'd87, 7'd55, 7'd31, 7'd59};
assign threshold_10[31] = 8'd56;
logic [4*types::LINE_BITS-1:0] line_11 [32];
logic [types::THRESH_BITS-1:0] threshold_11 [32];
assign line_11[0] = {7'd22, 7'd59, 7'd22, 7'd59};
assign threshold_11[0] = 8'd0;
assign line_11[1] = {7'd25, 7'd56, 7'd14, 7'd57};
assign threshold_11[1] = 8'd11;
assign line_11[2] = {7'd31, 7'd54, 7'd8, 7'd55};
assign threshold_11[2] = 8'd23;
assign line_11[3] = {7'd5, 7'd52, 7'd38, 7'd53};
assign threshold_11[3] = 8'd33;
assign line_11[4] = {7'd4, 7'd50, 7'd45, 7'd54};
assign threshold_11[4] = 8'd41;
assign line_11[5] = {7'd4, 7'd48, 7'd52, 7'd55};
assign threshold_11[5] = 8'd49;
assign line_11[6] = {7'd6, 7'd48, 7'd58, 7'd58};
assign threshold_11[6] = 8'd53;
assign line_11[7] = {7'd9, 7'd48, 7'd63, 7'd61};
assign threshold_11[7] = 8'd56;
assign line_11[8] = {7'd13, 7'd49, 7'd66, 7'd65};
assign threshold_11[8] = 8'd55;
assign line_11[9] = {7'd16, 7'd51, 7'd67, 7'd68};
assign threshold_11[9] = 8'd54;
assign line_11[10] = {7'd18, 7'd53, 7'd67, 7'd71};
assign threshold_11[10] = 8'd52;
assign line_11[11] = {7'd19, 7'd56, 7'd65, 7'd72};
assign threshold_11[11] = 8'd49;
assign line_11[12] = {7'd19, 7'd59, 7'd62, 7'd72};
assign threshold_11[12] = 8'd45;
assign line_11[13] = {7'd18, 7'd60, 7'd58, 7'd71};
assign threshold_11[13] = 8'd41;
assign line_11[14] = {7'd15, 7'd61, 7'd55, 7'd68};
assign threshold_11[14] = 8'd41;
assign line_11[15] = {7'd12, 7'd61, 7'd52, 7'd64};
assign threshold_11[15] = 8'd40;
assign line_11[16] = {7'd51, 7'd58, 7'd9, 7'd58};
assign threshold_11[16] = 8'd42;
assign line_11[17] = {7'd50, 7'd52, 7'd7, 7'd55};
assign threshold_11[17] = 8'd43;
assign line_11[18] = {7'd52, 7'd46, 7'd6, 7'd50};
assign threshold_11[18] = 8'd46;
assign line_11[19] = {7'd56, 7'd40, 7'd6, 7'd43};
assign threshold_11[19] = 8'd50;
assign line_11[20] = {7'd61, 7'd34, 7'd8, 7'd36};
assign threshold_11[20] = 8'd53;
assign line_11[21] = {7'd12, 7'd29, 7'd67, 7'd30};
assign threshold_11[21] = 8'd55;
assign line_11[22] = {7'd18, 7'd22, 7'd74, 7'd27};
assign threshold_11[22] = 8'd56;
assign line_11[23] = {7'd26, 7'd15, 7'd82, 7'd26};
assign threshold_11[23] = 8'd57;
assign line_11[24] = {7'd35, 7'd10, 7'd88, 7'd26};
assign threshold_11[24] = 8'd55;
assign line_11[25] = {7'd45, 7'd6, 7'd94, 7'd28};
assign threshold_11[25] = 8'd54;
assign line_11[26] = {7'd54, 7'd4, 7'd98, 7'd31};
assign threshold_11[26] = 8'd52;
assign line_11[27] = {7'd64, 7'd4, 7'd100, 7'd35};
assign threshold_11[27] = 8'd48;
assign line_11[28] = {7'd71, 7'd5, 7'd100, 7'd40};
assign threshold_11[28] = 8'd45;
assign line_11[29] = {7'd77, 7'd7, 7'd98, 7'd46};
assign threshold_11[29] = 8'd44;
assign line_11[30] = {7'd80, 7'd10, 7'd94, 7'd50};
assign threshold_11[30] = 8'd42;
assign line_11[31] = {7'd81, 7'd13, 7'd87, 7'd55};
assign threshold_11[31] = 8'd42;

endmodule
