// SPDX-FileCopyrightText: © 2024 Leo Moser <leo.moser@pm.me>
// SPDX-License-Identifier: Apache-2.0

`default_nettype none

module line_rom (
    input  logic [4:0] frame_i, // 32 frames
    input  logic [3:0] line_i,  // 12 lines
    
    output types::line_t      my_line,
    output logic [types::THRESH_BITS-1:0] my_thresh
);
    // Line
    always_comb begin
        case (line_i)
            4'd0: my_line = {point_0_x[frame_i], point_0_y[frame_i], point_1_x[frame_i], point_1_y[frame_i]};
            4'd1: my_line = {point_1_x[frame_i], point_1_y[frame_i], point_3_x[frame_i], point_3_y[frame_i]};
            4'd2: my_line = {point_3_x[frame_i], point_3_y[frame_i], point_2_x[frame_i], point_2_y[frame_i]};
            4'd3: my_line = {point_2_x[frame_i], point_2_y[frame_i], point_0_x[frame_i], point_0_y[frame_i]};
            4'd4: my_line = {point_0_x[frame_i], point_0_y[frame_i], point_4_x[frame_i], point_4_y[frame_i]};
            4'd5: my_line = {point_1_x[frame_i], point_1_y[frame_i], point_5_x[frame_i], point_5_y[frame_i]};
            4'd6: my_line = {point_2_x[frame_i], point_2_y[frame_i], point_6_x[frame_i], point_6_y[frame_i]};
            4'd7: my_line = {point_3_x[frame_i], point_3_y[frame_i], point_7_x[frame_i], point_7_y[frame_i]};
            4'd8: my_line = {point_4_x[frame_i], point_4_y[frame_i], point_5_x[frame_i], point_5_y[frame_i]};
            4'd9: my_line = {point_5_x[frame_i], point_5_y[frame_i], point_7_x[frame_i], point_7_y[frame_i]};
            4'd10: my_line = {point_7_x[frame_i], point_7_y[frame_i], point_6_x[frame_i], point_6_y[frame_i]};
            4'd11: my_line = {point_6_x[frame_i], point_6_y[frame_i], point_4_x[frame_i], point_4_y[frame_i]};
            default: my_line = 'x;
        endcase
    end
    
    // Threshold must be shifted because of the 
    // pipeline latency in the edge_function
    always_comb begin
        case (line_i)
            4'd0: my_thresh = threshold_10[frame_i];
            4'd1: my_thresh = threshold_11[frame_i];
            4'd2: my_thresh = threshold_0[frame_i];
            4'd3: my_thresh = threshold_1[frame_i];
            4'd4: my_thresh = threshold_2[frame_i];
            4'd5: my_thresh = threshold_3[frame_i];
            4'd6: my_thresh = threshold_4[frame_i];
            4'd7: my_thresh = threshold_5[frame_i];
            4'd8: my_thresh = threshold_6[frame_i];
            4'd9: my_thresh = threshold_7[frame_i];
            4'd10: my_thresh = threshold_8[frame_i];
            4'd11: my_thresh = threshold_9[frame_i];
            default: my_thresh = 'x;
        endcase
    end
    /*always_comb begin
        case (line_i)
            4'd0: my_thresh = threshold_9[frame_i];
            4'd1: my_thresh = threshold_10[frame_i];
            4'd2: my_thresh = threshold_11[frame_i];
            4'd3: my_thresh = threshold_0[frame_i];
            4'd4: my_thresh = threshold_1[frame_i];
            4'd5: my_thresh = threshold_2[frame_i];
            4'd6: my_thresh = threshold_3[frame_i];
            4'd7: my_thresh = threshold_4[frame_i];
            4'd8: my_thresh = threshold_5[frame_i];
            4'd9: my_thresh = threshold_6[frame_i];
            4'd10: my_thresh = threshold_7[frame_i];
            4'd11: my_thresh = threshold_8[frame_i];
            default: my_thresh = 'x;
        endcase
    end*/
    /*always_comb begin
        case (line_i)
            4'd0: my_thresh = threshold_8[frame_i];
            4'd1: my_thresh = threshold_9[frame_i];
            4'd2: my_thresh = threshold_10[frame_i];
            4'd3: my_thresh = threshold_11[frame_i];
            4'd4: my_thresh = threshold_0[frame_i];
            4'd5: my_thresh = threshold_1[frame_i];
            4'd6: my_thresh = threshold_2[frame_i];
            4'd7: my_thresh = threshold_3[frame_i];
            4'd8: my_thresh = threshold_4[frame_i];
            4'd9: my_thresh = threshold_5[frame_i];
            4'd10: my_thresh = threshold_6[frame_i];
            4'd11: my_thresh = threshold_7[frame_i];
            default: my_thresh = 'x;
        endcase
    end*/
    
logic [types::LINE_BITS-1:0] point_0_x [32];
logic [types::LINE_BITS-1:0] point_0_y [32];
assign point_0_x[0] = 7'd22;
assign point_0_y[0] = 7'd17;
assign point_0_x[1] = 7'd19;
assign point_0_y[1] = 7'd15;
assign point_0_x[2] = 7'd17;
assign point_0_y[2] = 7'd14;
assign point_0_x[3] = 7'd17;
assign point_0_y[3] = 7'd12;
assign point_0_x[4] = 7'd18;
assign point_0_y[4] = 7'd10;
assign point_0_x[5] = 7'd20;
assign point_0_y[5] = 7'd9;
assign point_0_x[6] = 7'd24;
assign point_0_y[6] = 7'd8;
assign point_0_x[7] = 7'd29;
assign point_0_y[7] = 7'd8;
assign point_0_x[8] = 7'd35;
assign point_0_y[8] = 7'd10;
assign point_0_x[9] = 7'd41;
assign point_0_y[9] = 7'd13;
assign point_0_x[10] = 7'd46;
assign point_0_y[10] = 7'd18;
assign point_0_x[11] = 7'd51;
assign point_0_y[11] = 7'd23;
assign point_0_x[12] = 7'd55;
assign point_0_y[12] = 7'd30;
assign point_0_x[13] = 7'd57;
assign point_0_y[13] = 7'd37;
assign point_0_x[14] = 7'd57;
assign point_0_y[14] = 7'd45;
assign point_0_x[15] = 7'd55;
assign point_0_y[15] = 7'd52;
assign point_0_x[16] = 7'd50;
assign point_0_y[16] = 7'd59;
assign point_0_x[17] = 7'd45;
assign point_0_y[17] = 7'd64;
assign point_0_x[18] = 7'd38;
assign point_0_y[18] = 7'd67;
assign point_0_x[19] = 7'd31;
assign point_0_y[19] = 7'd69;
assign point_0_x[20] = 7'd24;
assign point_0_y[20] = 7'd68;
assign point_0_x[21] = 7'd19;
assign point_0_y[21] = 7'd66;
assign point_0_x[22] = 7'd14;
assign point_0_y[22] = 7'd61;
assign point_0_x[23] = 7'd12;
assign point_0_y[23] = 7'd56;
assign point_0_x[24] = 7'd13;
assign point_0_y[24] = 7'd49;
assign point_0_x[25] = 7'd16;
assign point_0_y[25] = 7'd42;
assign point_0_x[26] = 7'd21;
assign point_0_y[26] = 7'd35;
assign point_0_x[27] = 7'd29;
assign point_0_y[27] = 7'd29;
assign point_0_x[28] = 7'd38;
assign point_0_y[28] = 7'd23;
assign point_0_x[29] = 7'd49;
assign point_0_y[29] = 7'd19;
assign point_0_x[30] = 7'd60;
assign point_0_y[30] = 7'd17;
assign point_0_x[31] = 7'd70;
assign point_0_y[31] = 7'd16;
logic [types::LINE_BITS-1:0] point_1_x [32];
logic [types::LINE_BITS-1:0] point_1_y [32];
assign point_1_x[0] = 7'd80;
assign point_1_y[0] = 7'd17;
assign point_1_x[1] = 7'd76;
assign point_1_y[1] = 7'd19;
assign point_1_x[2] = 7'd70;
assign point_1_y[2] = 7'd21;
assign point_1_x[3] = 7'd63;
assign point_1_y[3] = 7'd22;
assign point_1_x[4] = 7'd56;
assign point_1_y[4] = 7'd21;
assign point_1_x[5] = 7'd49;
assign point_1_y[5] = 7'd20;
assign point_1_x[6] = 7'd43;
assign point_1_y[6] = 7'd17;
assign point_1_x[7] = 7'd38;
assign point_1_y[7] = 7'd14;
assign point_1_x[8] = 7'd35;
assign point_1_y[8] = 7'd10;
assign point_1_x[9] = 7'd34;
assign point_1_y[9] = 7'd7;
assign point_1_x[10] = 7'd34;
assign point_1_y[10] = 7'd4;
assign point_1_x[11] = 7'd36;
assign point_1_y[11] = 7'd3;
assign point_1_x[12] = 7'd39;
assign point_1_y[12] = 7'd3;
assign point_1_x[13] = 7'd43;
assign point_1_y[13] = 7'd4;
assign point_1_x[14] = 7'd46;
assign point_1_y[14] = 7'd7;
assign point_1_x[15] = 7'd49;
assign point_1_y[15] = 7'd11;
assign point_1_x[16] = 7'd51;
assign point_1_y[16] = 7'd17;
assign point_1_x[17] = 7'd51;
assign point_1_y[17] = 7'd23;
assign point_1_x[18] = 7'd49;
assign point_1_y[18] = 7'd29;
assign point_1_x[19] = 7'd45;
assign point_1_y[19] = 7'd35;
assign point_1_x[20] = 7'd40;
assign point_1_y[20] = 7'd41;
assign point_1_x[21] = 7'd34;
assign point_1_y[21] = 7'd45;
assign point_1_x[22] = 7'd27;
assign point_1_y[22] = 7'd48;
assign point_1_x[23] = 7'd19;
assign point_1_y[23] = 7'd49;
assign point_1_x[24] = 7'd13;
assign point_1_y[24] = 7'd49;
assign point_1_x[25] = 7'd7;
assign point_1_y[25] = 7'd47;
assign point_1_x[26] = 7'd3;
assign point_1_y[26] = 7'd44;
assign point_1_x[27] = 7'd1;
assign point_1_y[27] = 7'd40;
assign point_1_x[28] = 7'd1;
assign point_1_y[28] = 7'd35;
assign point_1_x[29] = 7'd3;
assign point_1_y[29] = 7'd29;
assign point_1_x[30] = 7'd7;
assign point_1_y[30] = 7'd25;
assign point_1_x[31] = 7'd14;
assign point_1_y[31] = 7'd20;
logic [types::LINE_BITS-1:0] point_2_x [32];
logic [types::LINE_BITS-1:0] point_2_y [32];
assign point_2_x[0] = 7'd22;
assign point_2_y[0] = 7'd17;
assign point_2_x[1] = 7'd31;
assign point_2_y[1] = 7'd14;
assign point_2_x[2] = 7'd40;
assign point_2_y[2] = 7'd13;
assign point_2_x[3] = 7'd50;
assign point_2_y[3] = 7'd12;
assign point_2_x[4] = 7'd59;
assign point_2_y[4] = 7'd13;
assign point_2_x[5] = 7'd68;
assign point_2_y[5] = 7'd16;
assign point_2_x[6] = 7'd76;
assign point_2_y[6] = 7'd18;
assign point_2_x[7] = 7'd83;
assign point_2_y[7] = 7'd22;
assign point_2_x[8] = 7'd88;
assign point_2_y[8] = 7'd26;
assign point_2_x[9] = 7'd93;
assign point_2_y[9] = 7'd31;
assign point_2_x[10] = 7'd95;
assign point_2_y[10] = 7'd35;
assign point_2_x[11] = 7'd97;
assign point_2_y[11] = 7'd40;
assign point_2_x[12] = 7'd98;
assign point_2_y[12] = 7'd44;
assign point_2_x[13] = 7'd97;
assign point_2_y[13] = 7'd48;
assign point_2_x[14] = 7'd96;
assign point_2_y[14] = 7'd52;
assign point_2_x[15] = 7'd94;
assign point_2_y[15] = 7'd55;
assign point_2_x[16] = 7'd92;
assign point_2_y[16] = 7'd59;
assign point_2_x[17] = 7'd88;
assign point_2_y[17] = 7'd61;
assign point_2_x[18] = 7'd85;
assign point_2_y[18] = 7'd63;
assign point_2_x[19] = 7'd81;
assign point_2_y[19] = 7'd65;
assign point_2_x[20] = 7'd78;
assign point_2_y[20] = 7'd66;
assign point_2_x[21] = 7'd74;
assign point_2_y[21] = 7'd67;
assign point_2_x[22] = 7'd71;
assign point_2_y[22] = 7'd67;
assign point_2_x[23] = 7'd68;
assign point_2_y[23] = 7'd66;
assign point_2_x[24] = 7'd66;
assign point_2_y[24] = 7'd65;
assign point_2_x[25] = 7'd65;
assign point_2_y[25] = 7'd64;
assign point_2_x[26] = 7'd65;
assign point_2_y[26] = 7'd62;
assign point_2_x[27] = 7'd66;
assign point_2_y[27] = 7'd60;
assign point_2_x[28] = 7'd68;
assign point_2_y[28] = 7'd59;
assign point_2_x[29] = 7'd70;
assign point_2_y[29] = 7'd58;
assign point_2_x[30] = 7'd73;
assign point_2_y[30] = 7'd58;
assign point_2_x[31] = 7'd76;
assign point_2_y[31] = 7'd58;
logic [types::LINE_BITS-1:0] point_3_x [32];
logic [types::LINE_BITS-1:0] point_3_y [32];
assign point_3_x[0] = 7'd80;
assign point_3_y[0] = 7'd17;
assign point_3_x[1] = 7'd87;
assign point_3_y[1] = 7'd18;
assign point_3_x[2] = 7'd93;
assign point_3_y[2] = 7'd20;
assign point_3_x[3] = 7'd96;
assign point_3_y[3] = 7'd23;
assign point_3_x[4] = 7'd97;
assign point_3_y[4] = 7'd25;
assign point_3_x[5] = 7'd97;
assign point_3_y[5] = 7'd27;
assign point_3_x[6] = 7'd95;
assign point_3_y[6] = 7'd27;
assign point_3_x[7] = 7'd92;
assign point_3_y[7] = 7'd27;
assign point_3_x[8] = 7'd88;
assign point_3_y[8] = 7'd26;
assign point_3_x[9] = 7'd85;
assign point_3_y[9] = 7'd24;
assign point_3_x[10] = 7'd83;
assign point_3_y[10] = 7'd22;
assign point_3_x[11] = 7'd82;
assign point_3_y[11] = 7'd19;
assign point_3_x[12] = 7'd82;
assign point_3_y[12] = 7'd16;
assign point_3_x[13] = 7'd83;
assign point_3_y[13] = 7'd15;
assign point_3_x[14] = 7'd86;
assign point_3_y[14] = 7'd14;
assign point_3_x[15] = 7'd89;
assign point_3_y[15] = 7'd14;
assign point_3_x[16] = 7'd92;
assign point_3_y[16] = 7'd17;
assign point_3_x[17] = 7'd94;
assign point_3_y[17] = 7'd20;
assign point_3_x[18] = 7'd95;
assign point_3_y[18] = 7'd25;
assign point_3_x[19] = 7'd95;
assign point_3_y[19] = 7'd32;
assign point_3_x[20] = 7'd93;
assign point_3_y[20] = 7'd39;
assign point_3_x[21] = 7'd89;
assign point_3_y[21] = 7'd46;
assign point_3_x[22] = 7'd83;
assign point_3_y[22] = 7'd53;
assign point_3_x[23] = 7'd75;
assign point_3_y[23] = 7'd60;
assign point_3_x[24] = 7'd66;
assign point_3_y[24] = 7'd65;
assign point_3_x[25] = 7'd56;
assign point_3_y[25] = 7'd69;
assign point_3_x[26] = 7'd47;
assign point_3_y[26] = 7'd71;
assign point_3_x[27] = 7'd37;
assign point_3_y[27] = 7'd71;
assign point_3_x[28] = 7'd30;
assign point_3_y[28] = 7'd70;
assign point_3_x[29] = 7'd24;
assign point_3_y[29] = 7'd68;
assign point_3_x[30] = 7'd21;
assign point_3_y[30] = 7'd65;
assign point_3_x[31] = 7'd20;
assign point_3_y[31] = 7'd62;
logic [types::LINE_BITS-1:0] point_4_x [32];
logic [types::LINE_BITS-1:0] point_4_y [32];
assign point_4_x[0] = 7'd22;
assign point_4_y[0] = 7'd59;
assign point_4_x[1] = 7'd14;
assign point_4_y[1] = 7'd57;
assign point_4_x[2] = 7'd8;
assign point_4_y[2] = 7'd55;
assign point_4_x[3] = 7'd5;
assign point_4_y[3] = 7'd52;
assign point_4_x[4] = 7'd4;
assign point_4_y[4] = 7'd50;
assign point_4_x[5] = 7'd4;
assign point_4_y[5] = 7'd48;
assign point_4_x[6] = 7'd6;
assign point_4_y[6] = 7'd48;
assign point_4_x[7] = 7'd9;
assign point_4_y[7] = 7'd48;
assign point_4_x[8] = 7'd13;
assign point_4_y[8] = 7'd49;
assign point_4_x[9] = 7'd16;
assign point_4_y[9] = 7'd51;
assign point_4_x[10] = 7'd18;
assign point_4_y[10] = 7'd53;
assign point_4_x[11] = 7'd19;
assign point_4_y[11] = 7'd56;
assign point_4_x[12] = 7'd19;
assign point_4_y[12] = 7'd59;
assign point_4_x[13] = 7'd18;
assign point_4_y[13] = 7'd60;
assign point_4_x[14] = 7'd15;
assign point_4_y[14] = 7'd61;
assign point_4_x[15] = 7'd12;
assign point_4_y[15] = 7'd61;
assign point_4_x[16] = 7'd9;
assign point_4_y[16] = 7'd58;
assign point_4_x[17] = 7'd7;
assign point_4_y[17] = 7'd55;
assign point_4_x[18] = 7'd6;
assign point_4_y[18] = 7'd50;
assign point_4_x[19] = 7'd6;
assign point_4_y[19] = 7'd43;
assign point_4_x[20] = 7'd8;
assign point_4_y[20] = 7'd36;
assign point_4_x[21] = 7'd12;
assign point_4_y[21] = 7'd29;
assign point_4_x[22] = 7'd18;
assign point_4_y[22] = 7'd22;
assign point_4_x[23] = 7'd26;
assign point_4_y[23] = 7'd15;
assign point_4_x[24] = 7'd35;
assign point_4_y[24] = 7'd10;
assign point_4_x[25] = 7'd45;
assign point_4_y[25] = 7'd6;
assign point_4_x[26] = 7'd54;
assign point_4_y[26] = 7'd4;
assign point_4_x[27] = 7'd64;
assign point_4_y[27] = 7'd4;
assign point_4_x[28] = 7'd71;
assign point_4_y[28] = 7'd5;
assign point_4_x[29] = 7'd77;
assign point_4_y[29] = 7'd7;
assign point_4_x[30] = 7'd80;
assign point_4_y[30] = 7'd10;
assign point_4_x[31] = 7'd81;
assign point_4_y[31] = 7'd13;
logic [types::LINE_BITS-1:0] point_5_x [32];
logic [types::LINE_BITS-1:0] point_5_y [32];
assign point_5_x[0] = 7'd80;
assign point_5_y[0] = 7'd59;
assign point_5_x[1] = 7'd70;
assign point_5_y[1] = 7'd61;
assign point_5_x[2] = 7'd61;
assign point_5_y[2] = 7'd62;
assign point_5_x[3] = 7'd51;
assign point_5_y[3] = 7'd63;
assign point_5_x[4] = 7'd42;
assign point_5_y[4] = 7'd62;
assign point_5_x[5] = 7'd33;
assign point_5_y[5] = 7'd59;
assign point_5_x[6] = 7'd25;
assign point_5_y[6] = 7'd57;
assign point_5_x[7] = 7'd18;
assign point_5_y[7] = 7'd53;
assign point_5_x[8] = 7'd13;
assign point_5_y[8] = 7'd49;
assign point_5_x[9] = 7'd8;
assign point_5_y[9] = 7'd44;
assign point_5_x[10] = 7'd6;
assign point_5_y[10] = 7'd40;
assign point_5_x[11] = 7'd4;
assign point_5_y[11] = 7'd35;
assign point_5_x[12] = 7'd3;
assign point_5_y[12] = 7'd31;
assign point_5_x[13] = 7'd4;
assign point_5_y[13] = 7'd27;
assign point_5_x[14] = 7'd5;
assign point_5_y[14] = 7'd23;
assign point_5_x[15] = 7'd7;
assign point_5_y[15] = 7'd20;
assign point_5_x[16] = 7'd9;
assign point_5_y[16] = 7'd16;
assign point_5_x[17] = 7'd13;
assign point_5_y[17] = 7'd14;
assign point_5_x[18] = 7'd16;
assign point_5_y[18] = 7'd12;
assign point_5_x[19] = 7'd20;
assign point_5_y[19] = 7'd10;
assign point_5_x[20] = 7'd23;
assign point_5_y[20] = 7'd9;
assign point_5_x[21] = 7'd27;
assign point_5_y[21] = 7'd8;
assign point_5_x[22] = 7'd30;
assign point_5_y[22] = 7'd8;
assign point_5_x[23] = 7'd33;
assign point_5_y[23] = 7'd9;
assign point_5_x[24] = 7'd35;
assign point_5_y[24] = 7'd10;
assign point_5_x[25] = 7'd36;
assign point_5_y[25] = 7'd11;
assign point_5_x[26] = 7'd36;
assign point_5_y[26] = 7'd13;
assign point_5_x[27] = 7'd35;
assign point_5_y[27] = 7'd15;
assign point_5_x[28] = 7'd33;
assign point_5_y[28] = 7'd16;
assign point_5_x[29] = 7'd31;
assign point_5_y[29] = 7'd17;
assign point_5_x[30] = 7'd28;
assign point_5_y[30] = 7'd17;
assign point_5_x[31] = 7'd25;
assign point_5_y[31] = 7'd17;
logic [types::LINE_BITS-1:0] point_6_x [32];
logic [types::LINE_BITS-1:0] point_6_y [32];
assign point_6_x[0] = 7'd22;
assign point_6_y[0] = 7'd59;
assign point_6_x[1] = 7'd25;
assign point_6_y[1] = 7'd56;
assign point_6_x[2] = 7'd31;
assign point_6_y[2] = 7'd54;
assign point_6_x[3] = 7'd38;
assign point_6_y[3] = 7'd53;
assign point_6_x[4] = 7'd45;
assign point_6_y[4] = 7'd54;
assign point_6_x[5] = 7'd52;
assign point_6_y[5] = 7'd55;
assign point_6_x[6] = 7'd58;
assign point_6_y[6] = 7'd58;
assign point_6_x[7] = 7'd63;
assign point_6_y[7] = 7'd61;
assign point_6_x[8] = 7'd66;
assign point_6_y[8] = 7'd65;
assign point_6_x[9] = 7'd67;
assign point_6_y[9] = 7'd68;
assign point_6_x[10] = 7'd67;
assign point_6_y[10] = 7'd71;
assign point_6_x[11] = 7'd65;
assign point_6_y[11] = 7'd72;
assign point_6_x[12] = 7'd62;
assign point_6_y[12] = 7'd72;
assign point_6_x[13] = 7'd58;
assign point_6_y[13] = 7'd71;
assign point_6_x[14] = 7'd55;
assign point_6_y[14] = 7'd68;
assign point_6_x[15] = 7'd52;
assign point_6_y[15] = 7'd64;
assign point_6_x[16] = 7'd51;
assign point_6_y[16] = 7'd58;
assign point_6_x[17] = 7'd50;
assign point_6_y[17] = 7'd52;
assign point_6_x[18] = 7'd52;
assign point_6_y[18] = 7'd46;
assign point_6_x[19] = 7'd56;
assign point_6_y[19] = 7'd40;
assign point_6_x[20] = 7'd61;
assign point_6_y[20] = 7'd34;
assign point_6_x[21] = 7'd67;
assign point_6_y[21] = 7'd30;
assign point_6_x[22] = 7'd74;
assign point_6_y[22] = 7'd27;
assign point_6_x[23] = 7'd82;
assign point_6_y[23] = 7'd26;
assign point_6_x[24] = 7'd88;
assign point_6_y[24] = 7'd26;
assign point_6_x[25] = 7'd94;
assign point_6_y[25] = 7'd28;
assign point_6_x[26] = 7'd98;
assign point_6_y[26] = 7'd31;
assign point_6_x[27] = 7'd100;
assign point_6_y[27] = 7'd35;
assign point_6_x[28] = 7'd100;
assign point_6_y[28] = 7'd40;
assign point_6_x[29] = 7'd98;
assign point_6_y[29] = 7'd46;
assign point_6_x[30] = 7'd94;
assign point_6_y[30] = 7'd50;
assign point_6_x[31] = 7'd87;
assign point_6_y[31] = 7'd55;
logic [types::LINE_BITS-1:0] point_7_x [32];
logic [types::LINE_BITS-1:0] point_7_y [32];
assign point_7_x[0] = 7'd80;
assign point_7_y[0] = 7'd59;
assign point_7_x[1] = 7'd82;
assign point_7_y[1] = 7'd60;
assign point_7_x[2] = 7'd84;
assign point_7_y[2] = 7'd61;
assign point_7_x[3] = 7'd84;
assign point_7_y[3] = 7'd63;
assign point_7_x[4] = 7'd83;
assign point_7_y[4] = 7'd65;
assign point_7_x[5] = 7'd81;
assign point_7_y[5] = 7'd66;
assign point_7_x[6] = 7'd77;
assign point_7_y[6] = 7'd67;
assign point_7_x[7] = 7'd72;
assign point_7_y[7] = 7'd67;
assign point_7_x[8] = 7'd66;
assign point_7_y[8] = 7'd65;
assign point_7_x[9] = 7'd60;
assign point_7_y[9] = 7'd62;
assign point_7_x[10] = 7'd55;
assign point_7_y[10] = 7'd57;
assign point_7_x[11] = 7'd50;
assign point_7_y[11] = 7'd52;
assign point_7_x[12] = 7'd46;
assign point_7_y[12] = 7'd45;
assign point_7_x[13] = 7'd44;
assign point_7_y[13] = 7'd38;
assign point_7_x[14] = 7'd44;
assign point_7_y[14] = 7'd30;
assign point_7_x[15] = 7'd46;
assign point_7_y[15] = 7'd23;
assign point_7_x[16] = 7'd51;
assign point_7_y[16] = 7'd16;
assign point_7_x[17] = 7'd56;
assign point_7_y[17] = 7'd11;
assign point_7_x[18] = 7'd63;
assign point_7_y[18] = 7'd8;
assign point_7_x[19] = 7'd70;
assign point_7_y[19] = 7'd6;
assign point_7_x[20] = 7'd77;
assign point_7_y[20] = 7'd7;
assign point_7_x[21] = 7'd82;
assign point_7_y[21] = 7'd9;
assign point_7_x[22] = 7'd87;
assign point_7_y[22] = 7'd14;
assign point_7_x[23] = 7'd89;
assign point_7_y[23] = 7'd19;
assign point_7_x[24] = 7'd88;
assign point_7_y[24] = 7'd26;
assign point_7_x[25] = 7'd85;
assign point_7_y[25] = 7'd33;
assign point_7_x[26] = 7'd80;
assign point_7_y[26] = 7'd40;
assign point_7_x[27] = 7'd72;
assign point_7_y[27] = 7'd46;
assign point_7_x[28] = 7'd63;
assign point_7_y[28] = 7'd52;
assign point_7_x[29] = 7'd52;
assign point_7_y[29] = 7'd56;
assign point_7_x[30] = 7'd41;
assign point_7_y[30] = 7'd58;
assign point_7_x[31] = 7'd31;
assign point_7_y[31] = 7'd59;
logic [types::THRESH_BITS-1:0] threshold_0 [32];
assign threshold_0[0] = 8'd58;
assign threshold_0[1] = 8'd57;
assign threshold_0[2] = 8'd53;
assign threshold_0[3] = 8'd47;
assign threshold_0[4] = 8'd40;
assign threshold_0[5] = 8'd31;
assign threshold_0[6] = 8'd21;
assign threshold_0[7] = 8'd11;
assign threshold_0[8] = 8'd0;
assign threshold_0[9] = 8'd9;
assign threshold_0[10] = 8'd18;
assign threshold_0[11] = 8'd25;
assign threshold_0[12] = 8'd31;
assign threshold_0[13] = 8'd36;
assign threshold_0[14] = 8'd40;
assign threshold_0[15] = 8'd41;
assign threshold_0[16] = 8'd42;
assign threshold_0[17] = 8'd41;
assign threshold_0[18] = 8'd40;
assign threshold_0[19] = 8'd37;
assign threshold_0[20] = 8'd31;
assign threshold_0[21] = 8'd26;
assign threshold_0[22] = 8'd18;
assign threshold_0[23] = 8'd10;
assign threshold_0[24] = 8'd0;
assign threshold_0[25] = 8'd10;
assign threshold_0[26] = 8'd20;
assign threshold_0[27] = 8'd30;
assign threshold_0[28] = 8'd39;
assign threshold_0[29] = 8'd47;
assign threshold_0[30] = 8'd54;
assign threshold_0[31] = 8'd56;
logic [types::THRESH_BITS-1:0] threshold_1 [32];
assign threshold_1[0] = 8'd0;
assign threshold_1[1] = 8'd11;
assign threshold_1[2] = 8'd23;
assign threshold_1[3] = 8'd33;
assign threshold_1[4] = 8'd41;
assign threshold_1[5] = 8'd49;
assign threshold_1[6] = 8'd53;
assign threshold_1[7] = 8'd56;
assign threshold_1[8] = 8'd55;
assign threshold_1[9] = 8'd54;
assign threshold_1[10] = 8'd52;
assign threshold_1[11] = 8'd49;
assign threshold_1[12] = 8'd45;
assign threshold_1[13] = 8'd41;
assign threshold_1[14] = 8'd41;
assign threshold_1[15] = 8'd40;
assign threshold_1[16] = 8'd41;
assign threshold_1[17] = 8'd43;
assign threshold_1[18] = 8'd46;
assign threshold_1[19] = 8'd50;
assign threshold_1[20] = 8'd53;
assign threshold_1[21] = 8'd55;
assign threshold_1[22] = 8'd56;
assign threshold_1[23] = 8'd57;
assign threshold_1[24] = 8'd55;
assign threshold_1[25] = 8'd54;
assign threshold_1[26] = 8'd52;
assign threshold_1[27] = 8'd48;
assign threshold_1[28] = 8'd45;
assign threshold_1[29] = 8'd44;
assign threshold_1[30] = 8'd42;
assign threshold_1[31] = 8'd42;
logic [types::THRESH_BITS-1:0] threshold_2 [32];
assign threshold_2[0] = 8'd58;
assign threshold_2[1] = 8'd56;
assign threshold_2[2] = 8'd53;
assign threshold_2[3] = 8'd47;
assign threshold_2[4] = 8'd40;
assign threshold_2[5] = 8'd31;
assign threshold_2[6] = 8'd21;
assign threshold_2[7] = 8'd10;
assign threshold_2[8] = 8'd0;
assign threshold_2[9] = 8'd11;
assign threshold_2[10] = 8'd18;
assign threshold_2[11] = 8'd26;
assign threshold_2[12] = 8'd32;
assign threshold_2[13] = 8'd36;
assign threshold_2[14] = 8'd39;
assign threshold_2[15] = 8'd41;
assign threshold_2[16] = 8'd42;
assign threshold_2[17] = 8'd41;
assign threshold_2[18] = 8'd39;
assign threshold_2[19] = 8'd36;
assign threshold_2[20] = 8'd31;
assign threshold_2[21] = 8'd26;
assign threshold_2[22] = 8'd18;
assign threshold_2[23] = 8'd9;
assign threshold_2[24] = 8'd0;
assign threshold_2[25] = 8'd10;
assign threshold_2[26] = 8'd20;
assign threshold_2[27] = 8'd31;
assign threshold_2[28] = 8'd40;
assign threshold_2[29] = 8'd47;
assign threshold_2[30] = 8'd52;
assign threshold_2[31] = 8'd56;
logic [types::THRESH_BITS-1:0] threshold_3 [32];
assign threshold_3[0] = 8'd0;
assign threshold_3[1] = 8'd12;
assign threshold_3[2] = 8'd23;
assign threshold_3[3] = 8'd33;
assign threshold_3[4] = 8'd41;
assign threshold_3[5] = 8'd49;
assign threshold_3[6] = 8'd53;
assign threshold_3[7] = 8'd56;
assign threshold_3[8] = 8'd55;
assign threshold_3[9] = 8'd55;
assign threshold_3[10] = 8'd52;
assign threshold_3[11] = 8'd49;
assign threshold_3[12] = 8'd45;
assign threshold_3[13] = 8'd41;
assign threshold_3[14] = 8'd40;
assign threshold_3[15] = 8'd39;
assign threshold_3[16] = 8'd42;
assign threshold_3[17] = 8'd43;
assign threshold_3[18] = 8'd47;
assign threshold_3[19] = 8'd50;
assign threshold_3[20] = 8'd54;
assign threshold_3[21] = 8'd55;
assign threshold_3[22] = 8'd57;
assign threshold_3[23] = 8'd57;
assign threshold_3[24] = 8'd55;
assign threshold_3[25] = 8'd54;
assign threshold_3[26] = 8'd52;
assign threshold_3[27] = 8'd48;
assign threshold_3[28] = 8'd47;
assign threshold_3[29] = 8'd44;
assign threshold_3[30] = 8'd43;
assign threshold_3[31] = 8'd42;
logic [types::THRESH_BITS-1:0] threshold_4 [32];
assign threshold_4[0] = 8'd42;
assign threshold_4[1] = 8'd42;
assign threshold_4[2] = 8'd42;
assign threshold_4[3] = 8'd42;
assign threshold_4[4] = 8'd42;
assign threshold_4[5] = 8'd42;
assign threshold_4[6] = 8'd44;
assign threshold_4[7] = 8'd45;
assign threshold_4[8] = 8'd45;
assign threshold_4[9] = 8'd45;
assign threshold_4[10] = 8'd45;
assign threshold_4[11] = 8'd46;
assign threshold_4[12] = 8'd46;
assign threshold_4[13] = 8'd45;
assign threshold_4[14] = 8'd45;
assign threshold_4[15] = 8'd44;
assign threshold_4[16] = 8'd41;
assign threshold_4[17] = 8'd39;
assign threshold_4[18] = 8'd36;
assign threshold_4[19] = 8'd36;
assign threshold_4[20] = 8'd36;
assign threshold_4[21] = 8'd38;
assign threshold_4[22] = 8'd39;
assign threshold_4[23] = 8'd43;
assign threshold_4[24] = 8'd45;
assign threshold_4[25] = 8'd46;
assign threshold_4[26] = 8'd45;
assign threshold_4[27] = 8'd43;
assign threshold_4[28] = 8'd38;
assign threshold_4[29] = 8'd30;
assign threshold_4[30] = 8'd21;
assign threshold_4[31] = 8'd11;
logic [types::THRESH_BITS-1:0] threshold_5 [32];
assign threshold_5[0] = 8'd42;
assign threshold_5[1] = 8'd42;
assign threshold_5[2] = 8'd42;
assign threshold_5[3] = 8'd43;
assign threshold_5[4] = 8'd43;
assign threshold_5[5] = 8'd42;
assign threshold_5[6] = 8'd44;
assign threshold_5[7] = 8'd44;
assign threshold_5[8] = 8'd45;
assign threshold_5[9] = 8'd45;
assign threshold_5[10] = 8'd46;
assign threshold_5[11] = 8'd45;
assign threshold_5[12] = 8'd46;
assign threshold_5[13] = 8'd45;
assign threshold_5[14] = 8'd44;
assign threshold_5[15] = 8'd43;
assign threshold_5[16] = 8'd42;
assign threshold_5[17] = 8'd39;
assign threshold_5[18] = 8'd37;
assign threshold_5[19] = 8'd35;
assign threshold_5[20] = 8'd36;
assign threshold_5[21] = 8'd38;
assign threshold_5[22] = 8'd40;
assign threshold_5[23] = 8'd42;
assign threshold_5[24] = 8'd45;
assign threshold_5[25] = 8'd46;
assign threshold_5[26] = 8'd45;
assign threshold_5[27] = 8'd42;
assign threshold_5[28] = 8'd37;
assign threshold_5[29] = 8'd30;
assign threshold_5[30] = 8'd22;
assign threshold_5[31] = 8'd11;
logic [types::THRESH_BITS-1:0] threshold_6 [32];
assign threshold_6[0] = 8'd42;
assign threshold_6[1] = 8'd42;
assign threshold_6[2] = 8'd42;
assign threshold_6[3] = 8'd43;
assign threshold_6[4] = 8'd43;
assign threshold_6[5] = 8'd42;
assign threshold_6[6] = 8'd44;
assign threshold_6[7] = 8'd44;
assign threshold_6[8] = 8'd45;
assign threshold_6[9] = 8'd45;
assign threshold_6[10] = 8'd46;
assign threshold_6[11] = 8'd45;
assign threshold_6[12] = 8'd46;
assign threshold_6[13] = 8'd45;
assign threshold_6[14] = 8'd44;
assign threshold_6[15] = 8'd43;
assign threshold_6[16] = 8'd41;
assign threshold_6[17] = 8'd39;
assign threshold_6[18] = 8'd37;
assign threshold_6[19] = 8'd35;
assign threshold_6[20] = 8'd36;
assign threshold_6[21] = 8'd38;
assign threshold_6[22] = 8'd40;
assign threshold_6[23] = 8'd42;
assign threshold_6[24] = 8'd45;
assign threshold_6[25] = 8'd46;
assign threshold_6[26] = 8'd45;
assign threshold_6[27] = 8'd42;
assign threshold_6[28] = 8'd37;
assign threshold_6[29] = 8'd30;
assign threshold_6[30] = 8'd22;
assign threshold_6[31] = 8'd11;
logic [types::THRESH_BITS-1:0] threshold_7 [32];
assign threshold_7[0] = 8'd42;
assign threshold_7[1] = 8'd42;
assign threshold_7[2] = 8'd42;
assign threshold_7[3] = 8'd42;
assign threshold_7[4] = 8'd42;
assign threshold_7[5] = 8'd42;
assign threshold_7[6] = 8'd44;
assign threshold_7[7] = 8'd45;
assign threshold_7[8] = 8'd45;
assign threshold_7[9] = 8'd45;
assign threshold_7[10] = 8'd45;
assign threshold_7[11] = 8'd46;
assign threshold_7[12] = 8'd46;
assign threshold_7[13] = 8'd45;
assign threshold_7[14] = 8'd45;
assign threshold_7[15] = 8'd44;
assign threshold_7[16] = 8'd41;
assign threshold_7[17] = 8'd39;
assign threshold_7[18] = 8'd36;
assign threshold_7[19] = 8'd36;
assign threshold_7[20] = 8'd36;
assign threshold_7[21] = 8'd38;
assign threshold_7[22] = 8'd39;
assign threshold_7[23] = 8'd43;
assign threshold_7[24] = 8'd45;
assign threshold_7[25] = 8'd46;
assign threshold_7[26] = 8'd45;
assign threshold_7[27] = 8'd43;
assign threshold_7[28] = 8'd38;
assign threshold_7[29] = 8'd30;
assign threshold_7[30] = 8'd21;
assign threshold_7[31] = 8'd11;
logic [types::THRESH_BITS-1:0] threshold_8 [32];
assign threshold_8[0] = 8'd58;
assign threshold_8[1] = 8'd56;
assign threshold_8[2] = 8'd53;
assign threshold_8[3] = 8'd47;
assign threshold_8[4] = 8'd40;
assign threshold_8[5] = 8'd31;
assign threshold_8[6] = 8'd21;
assign threshold_8[7] = 8'd10;
assign threshold_8[8] = 8'd0;
assign threshold_8[9] = 8'd11;
assign threshold_8[10] = 8'd18;
assign threshold_8[11] = 8'd26;
assign threshold_8[12] = 8'd32;
assign threshold_8[13] = 8'd36;
assign threshold_8[14] = 8'd39;
assign threshold_8[15] = 8'd41;
assign threshold_8[16] = 8'd42;
assign threshold_8[17] = 8'd41;
assign threshold_8[18] = 8'd39;
assign threshold_8[19] = 8'd36;
assign threshold_8[20] = 8'd31;
assign threshold_8[21] = 8'd26;
assign threshold_8[22] = 8'd18;
assign threshold_8[23] = 8'd9;
assign threshold_8[24] = 8'd0;
assign threshold_8[25] = 8'd10;
assign threshold_8[26] = 8'd20;
assign threshold_8[27] = 8'd31;
assign threshold_8[28] = 8'd40;
assign threshold_8[29] = 8'd47;
assign threshold_8[30] = 8'd52;
assign threshold_8[31] = 8'd56;
logic [types::THRESH_BITS-1:0] threshold_9 [32];
assign threshold_9[0] = 8'd0;
assign threshold_9[1] = 8'd12;
assign threshold_9[2] = 8'd23;
assign threshold_9[3] = 8'd33;
assign threshold_9[4] = 8'd41;
assign threshold_9[5] = 8'd49;
assign threshold_9[6] = 8'd53;
assign threshold_9[7] = 8'd56;
assign threshold_9[8] = 8'd55;
assign threshold_9[9] = 8'd55;
assign threshold_9[10] = 8'd52;
assign threshold_9[11] = 8'd49;
assign threshold_9[12] = 8'd45;
assign threshold_9[13] = 8'd41;
assign threshold_9[14] = 8'd40;
assign threshold_9[15] = 8'd39;
assign threshold_9[16] = 8'd42;
assign threshold_9[17] = 8'd43;
assign threshold_9[18] = 8'd47;
assign threshold_9[19] = 8'd50;
assign threshold_9[20] = 8'd54;
assign threshold_9[21] = 8'd55;
assign threshold_9[22] = 8'd57;
assign threshold_9[23] = 8'd57;
assign threshold_9[24] = 8'd55;
assign threshold_9[25] = 8'd54;
assign threshold_9[26] = 8'd52;
assign threshold_9[27] = 8'd48;
assign threshold_9[28] = 8'd47;
assign threshold_9[29] = 8'd44;
assign threshold_9[30] = 8'd43;
assign threshold_9[31] = 8'd42;
logic [types::THRESH_BITS-1:0] threshold_10 [32];
assign threshold_10[0] = 8'd58;
assign threshold_10[1] = 8'd57;
assign threshold_10[2] = 8'd53;
assign threshold_10[3] = 8'd47;
assign threshold_10[4] = 8'd40;
assign threshold_10[5] = 8'd31;
assign threshold_10[6] = 8'd21;
assign threshold_10[7] = 8'd11;
assign threshold_10[8] = 8'd0;
assign threshold_10[9] = 8'd9;
assign threshold_10[10] = 8'd18;
assign threshold_10[11] = 8'd25;
assign threshold_10[12] = 8'd31;
assign threshold_10[13] = 8'd36;
assign threshold_10[14] = 8'd40;
assign threshold_10[15] = 8'd41;
assign threshold_10[16] = 8'd42;
assign threshold_10[17] = 8'd41;
assign threshold_10[18] = 8'd40;
assign threshold_10[19] = 8'd37;
assign threshold_10[20] = 8'd31;
assign threshold_10[21] = 8'd26;
assign threshold_10[22] = 8'd18;
assign threshold_10[23] = 8'd10;
assign threshold_10[24] = 8'd0;
assign threshold_10[25] = 8'd10;
assign threshold_10[26] = 8'd20;
assign threshold_10[27] = 8'd30;
assign threshold_10[28] = 8'd39;
assign threshold_10[29] = 8'd47;
assign threshold_10[30] = 8'd54;
assign threshold_10[31] = 8'd56;
logic [types::THRESH_BITS-1:0] threshold_11 [32];
assign threshold_11[0] = 8'd0;
assign threshold_11[1] = 8'd11;
assign threshold_11[2] = 8'd23;
assign threshold_11[3] = 8'd33;
assign threshold_11[4] = 8'd41;
assign threshold_11[5] = 8'd49;
assign threshold_11[6] = 8'd53;
assign threshold_11[7] = 8'd56;
assign threshold_11[8] = 8'd55;
assign threshold_11[9] = 8'd54;
assign threshold_11[10] = 8'd52;
assign threshold_11[11] = 8'd49;
assign threshold_11[12] = 8'd45;
assign threshold_11[13] = 8'd41;
assign threshold_11[14] = 8'd41;
assign threshold_11[15] = 8'd40;
assign threshold_11[16] = 8'd42;
assign threshold_11[17] = 8'd43;
assign threshold_11[18] = 8'd46;
assign threshold_11[19] = 8'd50;
assign threshold_11[20] = 8'd53;
assign threshold_11[21] = 8'd55;
assign threshold_11[22] = 8'd56;
assign threshold_11[23] = 8'd57;
assign threshold_11[24] = 8'd55;
assign threshold_11[25] = 8'd54;
assign threshold_11[26] = 8'd52;
assign threshold_11[27] = 8'd48;
assign threshold_11[28] = 8'd45;
assign threshold_11[29] = 8'd44;
assign threshold_11[30] = 8'd42;
assign threshold_11[31] = 8'd42;

endmodule
