// SPDX-FileCopyrightText: © 2024 Leo Moser <leo.moser@pm.me>
// SPDX-License-Identifier: Apache-2.0

`default_nettype none

module line_rom (
    input  logic [5:0] frame_i, // 64 frames
    input  logic [3:0] line_i,  // 12 lines
    
    output types::line_t      my_line,
    output logic [types::THRESH_BITS-1:0] my_thresh
);
    // Line
    always_comb begin
        case (line_i)
            4'd0: my_line = {point_0_x[frame_i], point_0_y[frame_i], point_1_x[frame_i], point_1_y[frame_i]};
            4'd1: my_line = {point_1_x[frame_i], point_1_y[frame_i], point_3_x[frame_i], point_3_y[frame_i]};
            4'd2: my_line = {point_3_x[frame_i], point_3_y[frame_i], point_2_x[frame_i], point_2_y[frame_i]};
            4'd3: my_line = {point_2_x[frame_i], point_2_y[frame_i], point_0_x[frame_i], point_0_y[frame_i]};
            4'd4: my_line = {point_0_x[frame_i], point_0_y[frame_i], point_4_x[frame_i], point_4_y[frame_i]};
            4'd5: my_line = {point_1_x[frame_i], point_1_y[frame_i], point_5_x[frame_i], point_5_y[frame_i]};
            4'd6: my_line = {point_2_x[frame_i], point_2_y[frame_i], point_6_x[frame_i], point_6_y[frame_i]};
            4'd7: my_line = {point_3_x[frame_i], point_3_y[frame_i], point_7_x[frame_i], point_7_y[frame_i]};
            4'd8: my_line = {point_4_x[frame_i], point_4_y[frame_i], point_5_x[frame_i], point_5_y[frame_i]};
            4'd9: my_line = {point_5_x[frame_i], point_5_y[frame_i], point_7_x[frame_i], point_7_y[frame_i]};
            4'd10: my_line = {point_7_x[frame_i], point_7_y[frame_i], point_6_x[frame_i], point_6_y[frame_i]};
            4'd11: my_line = {point_6_x[frame_i], point_6_y[frame_i], point_4_x[frame_i], point_4_y[frame_i]};
            default: my_line = 'x;
        endcase
    end
    
    // Threshold must be shifted because of the 
    // pipeline latency in the edge_function
    always_comb begin
        case (line_i)
            4'd0: my_thresh = threshold_9[frame_i];
            4'd1: my_thresh = threshold_10[frame_i];
            4'd2: my_thresh = threshold_11[frame_i];
            4'd3: my_thresh = threshold_0[frame_i];
            4'd4: my_thresh = threshold_1[frame_i];
            4'd5: my_thresh = threshold_2[frame_i];
            4'd6: my_thresh = threshold_3[frame_i];
            4'd7: my_thresh = threshold_4[frame_i];
            4'd8: my_thresh = threshold_5[frame_i];
            4'd9: my_thresh = threshold_6[frame_i];
            4'd10: my_thresh = threshold_7[frame_i];
            4'd11: my_thresh = threshold_8[frame_i];
            default: my_thresh = 'x;
        endcase
    end
    /*always_comb begin
        case (line_i)
            4'd0: my_thresh = threshold_8[frame_i];
            4'd1: my_thresh = threshold_9[frame_i];
            4'd2: my_thresh = threshold_10[frame_i];
            4'd3: my_thresh = threshold_11[frame_i];
            4'd4: my_thresh = threshold_0[frame_i];
            4'd5: my_thresh = threshold_1[frame_i];
            4'd6: my_thresh = threshold_2[frame_i];
            4'd7: my_thresh = threshold_3[frame_i];
            4'd8: my_thresh = threshold_4[frame_i];
            4'd9: my_thresh = threshold_5[frame_i];
            4'd10: my_thresh = threshold_6[frame_i];
            4'd11: my_thresh = threshold_7[frame_i];
            default: my_thresh = 'x;
        endcase
    end*/
    
logic [types::LINE_BITS-1:0] point_0_x [64];
logic [types::LINE_BITS-1:0] point_0_y [64];
assign point_0_x[0] = 7'd22;
assign point_0_y[0] = 7'd17;
assign point_0_x[1] = 7'd20;
assign point_0_y[1] = 7'd16;
assign point_0_x[2] = 7'd19;
assign point_0_y[2] = 7'd15;
assign point_0_x[3] = 7'd18;
assign point_0_y[3] = 7'd14;
assign point_0_x[4] = 7'd17;
assign point_0_y[4] = 7'd14;
assign point_0_x[5] = 7'd17;
assign point_0_y[5] = 7'd13;
assign point_0_x[6] = 7'd17;
assign point_0_y[6] = 7'd12;
assign point_0_x[7] = 7'd17;
assign point_0_y[7] = 7'd11;
assign point_0_x[8] = 7'd18;
assign point_0_y[8] = 7'd10;
assign point_0_x[9] = 7'd19;
assign point_0_y[9] = 7'd9;
assign point_0_x[10] = 7'd20;
assign point_0_y[10] = 7'd9;
assign point_0_x[11] = 7'd22;
assign point_0_y[11] = 7'd8;
assign point_0_x[12] = 7'd24;
assign point_0_y[12] = 7'd8;
assign point_0_x[13] = 7'd27;
assign point_0_y[13] = 7'd8;
assign point_0_x[14] = 7'd29;
assign point_0_y[14] = 7'd8;
assign point_0_x[15] = 7'd32;
assign point_0_y[15] = 7'd9;
assign point_0_x[16] = 7'd35;
assign point_0_y[16] = 7'd10;
assign point_0_x[17] = 7'd38;
assign point_0_y[17] = 7'd11;
assign point_0_x[18] = 7'd41;
assign point_0_y[18] = 7'd13;
assign point_0_x[19] = 7'd44;
assign point_0_y[19] = 7'd15;
assign point_0_x[20] = 7'd46;
assign point_0_y[20] = 7'd18;
assign point_0_x[21] = 7'd49;
assign point_0_y[21] = 7'd20;
assign point_0_x[22] = 7'd51;
assign point_0_y[22] = 7'd23;
assign point_0_x[23] = 7'd53;
assign point_0_y[23] = 7'd27;
assign point_0_x[24] = 7'd55;
assign point_0_y[24] = 7'd30;
assign point_0_x[25] = 7'd56;
assign point_0_y[25] = 7'd34;
assign point_0_x[26] = 7'd57;
assign point_0_y[26] = 7'd37;
assign point_0_x[27] = 7'd57;
assign point_0_y[27] = 7'd41;
assign point_0_x[28] = 7'd57;
assign point_0_y[28] = 7'd45;
assign point_0_x[29] = 7'd56;
assign point_0_y[29] = 7'd49;
assign point_0_x[30] = 7'd55;
assign point_0_y[30] = 7'd52;
assign point_0_x[31] = 7'd53;
assign point_0_y[31] = 7'd55;
assign point_0_x[32] = 7'd50;
assign point_0_y[32] = 7'd59;
assign point_0_x[33] = 7'd48;
assign point_0_y[33] = 7'd61;
assign point_0_x[34] = 7'd45;
assign point_0_y[34] = 7'd64;
assign point_0_x[35] = 7'd42;
assign point_0_y[35] = 7'd66;
assign point_0_x[36] = 7'd38;
assign point_0_y[36] = 7'd67;
assign point_0_x[37] = 7'd35;
assign point_0_y[37] = 7'd68;
assign point_0_x[38] = 7'd31;
assign point_0_y[38] = 7'd69;
assign point_0_x[39] = 7'd28;
assign point_0_y[39] = 7'd69;
assign point_0_x[40] = 7'd24;
assign point_0_y[40] = 7'd68;
assign point_0_x[41] = 7'd21;
assign point_0_y[41] = 7'd67;
assign point_0_x[42] = 7'd19;
assign point_0_y[42] = 7'd66;
assign point_0_x[43] = 7'd16;
assign point_0_y[43] = 7'd64;
assign point_0_x[44] = 7'd14;
assign point_0_y[44] = 7'd61;
assign point_0_x[45] = 7'd13;
assign point_0_y[45] = 7'd59;
assign point_0_x[46] = 7'd12;
assign point_0_y[46] = 7'd56;
assign point_0_x[47] = 7'd12;
assign point_0_y[47] = 7'd52;
assign point_0_x[48] = 7'd13;
assign point_0_y[48] = 7'd49;
assign point_0_x[49] = 7'd14;
assign point_0_y[49] = 7'd45;
assign point_0_x[50] = 7'd16;
assign point_0_y[50] = 7'd42;
assign point_0_x[51] = 7'd18;
assign point_0_y[51] = 7'd38;
assign point_0_x[52] = 7'd21;
assign point_0_y[52] = 7'd35;
assign point_0_x[53] = 7'd25;
assign point_0_y[53] = 7'd32;
assign point_0_x[54] = 7'd29;
assign point_0_y[54] = 7'd29;
assign point_0_x[55] = 7'd34;
assign point_0_y[55] = 7'd26;
assign point_0_x[56] = 7'd38;
assign point_0_y[56] = 7'd23;
assign point_0_x[57] = 7'd44;
assign point_0_y[57] = 7'd21;
assign point_0_x[58] = 7'd49;
assign point_0_y[58] = 7'd19;
assign point_0_x[59] = 7'd54;
assign point_0_y[59] = 7'd18;
assign point_0_x[60] = 7'd60;
assign point_0_y[60] = 7'd17;
assign point_0_x[61] = 7'd65;
assign point_0_y[61] = 7'd16;
assign point_0_x[62] = 7'd70;
assign point_0_y[62] = 7'd16;
assign point_0_x[63] = 7'd75;
assign point_0_y[63] = 7'd16;
logic [types::LINE_BITS-1:0] point_1_x [64];
logic [types::LINE_BITS-1:0] point_1_y [64];
assign point_1_x[0] = 7'd80;
assign point_1_y[0] = 7'd17;
assign point_1_x[1] = 7'd78;
assign point_1_y[1] = 7'd18;
assign point_1_x[2] = 7'd76;
assign point_1_y[2] = 7'd19;
assign point_1_x[3] = 7'd73;
assign point_1_y[3] = 7'd20;
assign point_1_x[4] = 7'd70;
assign point_1_y[4] = 7'd21;
assign point_1_x[5] = 7'd67;
assign point_1_y[5] = 7'd22;
assign point_1_x[6] = 7'd63;
assign point_1_y[6] = 7'd22;
assign point_1_x[7] = 7'd60;
assign point_1_y[7] = 7'd22;
assign point_1_x[8] = 7'd56;
assign point_1_y[8] = 7'd21;
assign point_1_x[9] = 7'd52;
assign point_1_y[9] = 7'd21;
assign point_1_x[10] = 7'd49;
assign point_1_y[10] = 7'd20;
assign point_1_x[11] = 7'd46;
assign point_1_y[11] = 7'd18;
assign point_1_x[12] = 7'd43;
assign point_1_y[12] = 7'd17;
assign point_1_x[13] = 7'd40;
assign point_1_y[13] = 7'd15;
assign point_1_x[14] = 7'd38;
assign point_1_y[14] = 7'd14;
assign point_1_x[15] = 7'd36;
assign point_1_y[15] = 7'd12;
assign point_1_x[16] = 7'd35;
assign point_1_y[16] = 7'd10;
assign point_1_x[17] = 7'd34;
assign point_1_y[17] = 7'd8;
assign point_1_x[18] = 7'd34;
assign point_1_y[18] = 7'd7;
assign point_1_x[19] = 7'd34;
assign point_1_y[19] = 7'd5;
assign point_1_x[20] = 7'd34;
assign point_1_y[20] = 7'd4;
assign point_1_x[21] = 7'd35;
assign point_1_y[21] = 7'd3;
assign point_1_x[22] = 7'd36;
assign point_1_y[22] = 7'd3;
assign point_1_x[23] = 7'd38;
assign point_1_y[23] = 7'd2;
assign point_1_x[24] = 7'd39;
assign point_1_y[24] = 7'd3;
assign point_1_x[25] = 7'd41;
assign point_1_y[25] = 7'd3;
assign point_1_x[26] = 7'd43;
assign point_1_y[26] = 7'd4;
assign point_1_x[27] = 7'd44;
assign point_1_y[27] = 7'd5;
assign point_1_x[28] = 7'd46;
assign point_1_y[28] = 7'd7;
assign point_1_x[29] = 7'd48;
assign point_1_y[29] = 7'd9;
assign point_1_x[30] = 7'd49;
assign point_1_y[30] = 7'd11;
assign point_1_x[31] = 7'd50;
assign point_1_y[31] = 7'd14;
assign point_1_x[32] = 7'd51;
assign point_1_y[32] = 7'd17;
assign point_1_x[33] = 7'd51;
assign point_1_y[33] = 7'd19;
assign point_1_x[34] = 7'd51;
assign point_1_y[34] = 7'd23;
assign point_1_x[35] = 7'd50;
assign point_1_y[35] = 7'd26;
assign point_1_x[36] = 7'd49;
assign point_1_y[36] = 7'd29;
assign point_1_x[37] = 7'd47;
assign point_1_y[37] = 7'd32;
assign point_1_x[38] = 7'd45;
assign point_1_y[38] = 7'd35;
assign point_1_x[39] = 7'd43;
assign point_1_y[39] = 7'd38;
assign point_1_x[40] = 7'd40;
assign point_1_y[40] = 7'd41;
assign point_1_x[41] = 7'd37;
assign point_1_y[41] = 7'd43;
assign point_1_x[42] = 7'd34;
assign point_1_y[42] = 7'd45;
assign point_1_x[43] = 7'd30;
assign point_1_y[43] = 7'd47;
assign point_1_x[44] = 7'd27;
assign point_1_y[44] = 7'd48;
assign point_1_x[45] = 7'd23;
assign point_1_y[45] = 7'd49;
assign point_1_x[46] = 7'd19;
assign point_1_y[46] = 7'd49;
assign point_1_x[47] = 7'd16;
assign point_1_y[47] = 7'd49;
assign point_1_x[48] = 7'd13;
assign point_1_y[48] = 7'd49;
assign point_1_x[49] = 7'd10;
assign point_1_y[49] = 7'd48;
assign point_1_x[50] = 7'd7;
assign point_1_y[50] = 7'd47;
assign point_1_x[51] = 7'd5;
assign point_1_y[51] = 7'd46;
assign point_1_x[52] = 7'd3;
assign point_1_y[52] = 7'd44;
assign point_1_x[53] = 7'd1;
assign point_1_y[53] = 7'd42;
assign point_1_x[54] = 7'd1;
assign point_1_y[54] = 7'd40;
assign point_1_x[55] = 7'd0;
assign point_1_y[55] = 7'd37;
assign point_1_x[56] = 7'd1;
assign point_1_y[56] = 7'd35;
assign point_1_x[57] = 7'd1;
assign point_1_y[57] = 7'd32;
assign point_1_x[58] = 7'd3;
assign point_1_y[58] = 7'd29;
assign point_1_x[59] = 7'd5;
assign point_1_y[59] = 7'd27;
assign point_1_x[60] = 7'd7;
assign point_1_y[60] = 7'd25;
assign point_1_x[61] = 7'd10;
assign point_1_y[61] = 7'd22;
assign point_1_x[62] = 7'd14;
assign point_1_y[62] = 7'd20;
assign point_1_x[63] = 7'd17;
assign point_1_y[63] = 7'd18;
logic [types::LINE_BITS-1:0] point_2_x [64];
logic [types::LINE_BITS-1:0] point_2_y [64];
assign point_2_x[0] = 7'd22;
assign point_2_y[0] = 7'd17;
assign point_2_x[1] = 7'd26;
assign point_2_y[1] = 7'd15;
assign point_2_x[2] = 7'd31;
assign point_2_y[2] = 7'd14;
assign point_2_x[3] = 7'd35;
assign point_2_y[3] = 7'd13;
assign point_2_x[4] = 7'd40;
assign point_2_y[4] = 7'd13;
assign point_2_x[5] = 7'd45;
assign point_2_y[5] = 7'd12;
assign point_2_x[6] = 7'd50;
assign point_2_y[6] = 7'd12;
assign point_2_x[7] = 7'd55;
assign point_2_y[7] = 7'd13;
assign point_2_x[8] = 7'd59;
assign point_2_y[8] = 7'd13;
assign point_2_x[9] = 7'd64;
assign point_2_y[9] = 7'd14;
assign point_2_x[10] = 7'd68;
assign point_2_y[10] = 7'd16;
assign point_2_x[11] = 7'd72;
assign point_2_y[11] = 7'd17;
assign point_2_x[12] = 7'd76;
assign point_2_y[12] = 7'd18;
assign point_2_x[13] = 7'd80;
assign point_2_y[13] = 7'd20;
assign point_2_x[14] = 7'd83;
assign point_2_y[14] = 7'd22;
assign point_2_x[15] = 7'd86;
assign point_2_y[15] = 7'd24;
assign point_2_x[16] = 7'd88;
assign point_2_y[16] = 7'd26;
assign point_2_x[17] = 7'd91;
assign point_2_y[17] = 7'd28;
assign point_2_x[18] = 7'd93;
assign point_2_y[18] = 7'd31;
assign point_2_x[19] = 7'd94;
assign point_2_y[19] = 7'd33;
assign point_2_x[20] = 7'd95;
assign point_2_y[20] = 7'd35;
assign point_2_x[21] = 7'd96;
assign point_2_y[21] = 7'd37;
assign point_2_x[22] = 7'd97;
assign point_2_y[22] = 7'd40;
assign point_2_x[23] = 7'd98;
assign point_2_y[23] = 7'd42;
assign point_2_x[24] = 7'd98;
assign point_2_y[24] = 7'd44;
assign point_2_x[25] = 7'd98;
assign point_2_y[25] = 7'd46;
assign point_2_x[26] = 7'd97;
assign point_2_y[26] = 7'd48;
assign point_2_x[27] = 7'd97;
assign point_2_y[27] = 7'd50;
assign point_2_x[28] = 7'd96;
assign point_2_y[28] = 7'd52;
assign point_2_x[29] = 7'd95;
assign point_2_y[29] = 7'd54;
assign point_2_x[30] = 7'd94;
assign point_2_y[30] = 7'd55;
assign point_2_x[31] = 7'd93;
assign point_2_y[31] = 7'd57;
assign point_2_x[32] = 7'd92;
assign point_2_y[32] = 7'd59;
assign point_2_x[33] = 7'd90;
assign point_2_y[33] = 7'd60;
assign point_2_x[34] = 7'd88;
assign point_2_y[34] = 7'd61;
assign point_2_x[35] = 7'd87;
assign point_2_y[35] = 7'd62;
assign point_2_x[36] = 7'd85;
assign point_2_y[36] = 7'd63;
assign point_2_x[37] = 7'd83;
assign point_2_y[37] = 7'd64;
assign point_2_x[38] = 7'd81;
assign point_2_y[38] = 7'd65;
assign point_2_x[39] = 7'd79;
assign point_2_y[39] = 7'd66;
assign point_2_x[40] = 7'd78;
assign point_2_y[40] = 7'd66;
assign point_2_x[41] = 7'd76;
assign point_2_y[41] = 7'd66;
assign point_2_x[42] = 7'd74;
assign point_2_y[42] = 7'd67;
assign point_2_x[43] = 7'd72;
assign point_2_y[43] = 7'd67;
assign point_2_x[44] = 7'd71;
assign point_2_y[44] = 7'd67;
assign point_2_x[45] = 7'd69;
assign point_2_y[45] = 7'd66;
assign point_2_x[46] = 7'd68;
assign point_2_y[46] = 7'd66;
assign point_2_x[47] = 7'd67;
assign point_2_y[47] = 7'd66;
assign point_2_x[48] = 7'd66;
assign point_2_y[48] = 7'd65;
assign point_2_x[49] = 7'd66;
assign point_2_y[49] = 7'd64;
assign point_2_x[50] = 7'd65;
assign point_2_y[50] = 7'd64;
assign point_2_x[51] = 7'd65;
assign point_2_y[51] = 7'd63;
assign point_2_x[52] = 7'd65;
assign point_2_y[52] = 7'd62;
assign point_2_x[53] = 7'd65;
assign point_2_y[53] = 7'd61;
assign point_2_x[54] = 7'd66;
assign point_2_y[54] = 7'd60;
assign point_2_x[55] = 7'd67;
assign point_2_y[55] = 7'd60;
assign point_2_x[56] = 7'd68;
assign point_2_y[56] = 7'd59;
assign point_2_x[57] = 7'd69;
assign point_2_y[57] = 7'd59;
assign point_2_x[58] = 7'd70;
assign point_2_y[58] = 7'd58;
assign point_2_x[59] = 7'd72;
assign point_2_y[59] = 7'd58;
assign point_2_x[60] = 7'd73;
assign point_2_y[60] = 7'd58;
assign point_2_x[61] = 7'd75;
assign point_2_y[61] = 7'd58;
assign point_2_x[62] = 7'd76;
assign point_2_y[62] = 7'd58;
assign point_2_x[63] = 7'd78;
assign point_2_y[63] = 7'd58;
logic [types::LINE_BITS-1:0] point_3_x [64];
logic [types::LINE_BITS-1:0] point_3_y [64];
assign point_3_x[0] = 7'd80;
assign point_3_y[0] = 7'd17;
assign point_3_x[1] = 7'd84;
assign point_3_y[1] = 7'd17;
assign point_3_x[2] = 7'd87;
assign point_3_y[2] = 7'd18;
assign point_3_x[3] = 7'd90;
assign point_3_y[3] = 7'd19;
assign point_3_x[4] = 7'd93;
assign point_3_y[4] = 7'd20;
assign point_3_x[5] = 7'd95;
assign point_3_y[5] = 7'd21;
assign point_3_x[6] = 7'd96;
assign point_3_y[6] = 7'd23;
assign point_3_x[7] = 7'd97;
assign point_3_y[7] = 7'd24;
assign point_3_x[8] = 7'd97;
assign point_3_y[8] = 7'd25;
assign point_3_x[9] = 7'd97;
assign point_3_y[9] = 7'd26;
assign point_3_x[10] = 7'd97;
assign point_3_y[10] = 7'd27;
assign point_3_x[11] = 7'd96;
assign point_3_y[11] = 7'd27;
assign point_3_x[12] = 7'd95;
assign point_3_y[12] = 7'd27;
assign point_3_x[13] = 7'd93;
assign point_3_y[13] = 7'd27;
assign point_3_x[14] = 7'd92;
assign point_3_y[14] = 7'd27;
assign point_3_x[15] = 7'd90;
assign point_3_y[15] = 7'd27;
assign point_3_x[16] = 7'd88;
assign point_3_y[16] = 7'd26;
assign point_3_x[17] = 7'd87;
assign point_3_y[17] = 7'd25;
assign point_3_x[18] = 7'd85;
assign point_3_y[18] = 7'd24;
assign point_3_x[19] = 7'd84;
assign point_3_y[19] = 7'd23;
assign point_3_x[20] = 7'd83;
assign point_3_y[20] = 7'd22;
assign point_3_x[21] = 7'd82;
assign point_3_y[21] = 7'd20;
assign point_3_x[22] = 7'd82;
assign point_3_y[22] = 7'd19;
assign point_3_x[23] = 7'd82;
assign point_3_y[23] = 7'd18;
assign point_3_x[24] = 7'd82;
assign point_3_y[24] = 7'd16;
assign point_3_x[25] = 7'd82;
assign point_3_y[25] = 7'd15;
assign point_3_x[26] = 7'd83;
assign point_3_y[26] = 7'd15;
assign point_3_x[27] = 7'd84;
assign point_3_y[27] = 7'd14;
assign point_3_x[28] = 7'd86;
assign point_3_y[28] = 7'd14;
assign point_3_x[29] = 7'd87;
assign point_3_y[29] = 7'd14;
assign point_3_x[30] = 7'd89;
assign point_3_y[30] = 7'd14;
assign point_3_x[31] = 7'd90;
assign point_3_y[31] = 7'd15;
assign point_3_x[32] = 7'd92;
assign point_3_y[32] = 7'd17;
assign point_3_x[33] = 7'd93;
assign point_3_y[33] = 7'd18;
assign point_3_x[34] = 7'd94;
assign point_3_y[34] = 7'd20;
assign point_3_x[35] = 7'd95;
assign point_3_y[35] = 7'd23;
assign point_3_x[36] = 7'd95;
assign point_3_y[36] = 7'd25;
assign point_3_x[37] = 7'd96;
assign point_3_y[37] = 7'd28;
assign point_3_x[38] = 7'd95;
assign point_3_y[38] = 7'd32;
assign point_3_x[39] = 7'd95;
assign point_3_y[39] = 7'd35;
assign point_3_x[40] = 7'd93;
assign point_3_y[40] = 7'd39;
assign point_3_x[41] = 7'd92;
assign point_3_y[41] = 7'd42;
assign point_3_x[42] = 7'd89;
assign point_3_y[42] = 7'd46;
assign point_3_x[43] = 7'd86;
assign point_3_y[43] = 7'd50;
assign point_3_x[44] = 7'd83;
assign point_3_y[44] = 7'd53;
assign point_3_x[45] = 7'd79;
assign point_3_y[45] = 7'd57;
assign point_3_x[46] = 7'd75;
assign point_3_y[46] = 7'd60;
assign point_3_x[47] = 7'd71;
assign point_3_y[47] = 7'd62;
assign point_3_x[48] = 7'd66;
assign point_3_y[48] = 7'd65;
assign point_3_x[49] = 7'd61;
assign point_3_y[49] = 7'd67;
assign point_3_x[50] = 7'd56;
assign point_3_y[50] = 7'd69;
assign point_3_x[51] = 7'd51;
assign point_3_y[51] = 7'd70;
assign point_3_x[52] = 7'd47;
assign point_3_y[52] = 7'd71;
assign point_3_x[53] = 7'd42;
assign point_3_y[53] = 7'd71;
assign point_3_x[54] = 7'd37;
assign point_3_y[54] = 7'd71;
assign point_3_x[55] = 7'd33;
assign point_3_y[55] = 7'd71;
assign point_3_x[56] = 7'd30;
assign point_3_y[56] = 7'd70;
assign point_3_x[57] = 7'd27;
assign point_3_y[57] = 7'd69;
assign point_3_x[58] = 7'd24;
assign point_3_y[58] = 7'd68;
assign point_3_x[59] = 7'd22;
assign point_3_y[59] = 7'd67;
assign point_3_x[60] = 7'd21;
assign point_3_y[60] = 7'd65;
assign point_3_x[61] = 7'd20;
assign point_3_y[61] = 7'd64;
assign point_3_x[62] = 7'd20;
assign point_3_y[62] = 7'd62;
assign point_3_x[63] = 7'd20;
assign point_3_y[63] = 7'd60;
logic [types::LINE_BITS-1:0] point_4_x [64];
logic [types::LINE_BITS-1:0] point_4_y [64];
assign point_4_x[0] = 7'd22;
assign point_4_y[0] = 7'd59;
assign point_4_x[1] = 7'd17;
assign point_4_y[1] = 7'd58;
assign point_4_x[2] = 7'd14;
assign point_4_y[2] = 7'd57;
assign point_4_x[3] = 7'd11;
assign point_4_y[3] = 7'd56;
assign point_4_x[4] = 7'd8;
assign point_4_y[4] = 7'd55;
assign point_4_x[5] = 7'd6;
assign point_4_y[5] = 7'd54;
assign point_4_x[6] = 7'd5;
assign point_4_y[6] = 7'd52;
assign point_4_x[7] = 7'd4;
assign point_4_y[7] = 7'd51;
assign point_4_x[8] = 7'd4;
assign point_4_y[8] = 7'd50;
assign point_4_x[9] = 7'd4;
assign point_4_y[9] = 7'd49;
assign point_4_x[10] = 7'd4;
assign point_4_y[10] = 7'd48;
assign point_4_x[11] = 7'd5;
assign point_4_y[11] = 7'd48;
assign point_4_x[12] = 7'd6;
assign point_4_y[12] = 7'd48;
assign point_4_x[13] = 7'd8;
assign point_4_y[13] = 7'd48;
assign point_4_x[14] = 7'd9;
assign point_4_y[14] = 7'd48;
assign point_4_x[15] = 7'd11;
assign point_4_y[15] = 7'd48;
assign point_4_x[16] = 7'd13;
assign point_4_y[16] = 7'd49;
assign point_4_x[17] = 7'd14;
assign point_4_y[17] = 7'd50;
assign point_4_x[18] = 7'd16;
assign point_4_y[18] = 7'd51;
assign point_4_x[19] = 7'd17;
assign point_4_y[19] = 7'd52;
assign point_4_x[20] = 7'd18;
assign point_4_y[20] = 7'd53;
assign point_4_x[21] = 7'd19;
assign point_4_y[21] = 7'd55;
assign point_4_x[22] = 7'd19;
assign point_4_y[22] = 7'd56;
assign point_4_x[23] = 7'd19;
assign point_4_y[23] = 7'd57;
assign point_4_x[24] = 7'd19;
assign point_4_y[24] = 7'd59;
assign point_4_x[25] = 7'd19;
assign point_4_y[25] = 7'd60;
assign point_4_x[26] = 7'd18;
assign point_4_y[26] = 7'd60;
assign point_4_x[27] = 7'd17;
assign point_4_y[27] = 7'd61;
assign point_4_x[28] = 7'd15;
assign point_4_y[28] = 7'd61;
assign point_4_x[29] = 7'd14;
assign point_4_y[29] = 7'd61;
assign point_4_x[30] = 7'd12;
assign point_4_y[30] = 7'd61;
assign point_4_x[31] = 7'd11;
assign point_4_y[31] = 7'd60;
assign point_4_x[32] = 7'd9;
assign point_4_y[32] = 7'd58;
assign point_4_x[33] = 7'd8;
assign point_4_y[33] = 7'd57;
assign point_4_x[34] = 7'd7;
assign point_4_y[34] = 7'd55;
assign point_4_x[35] = 7'd6;
assign point_4_y[35] = 7'd52;
assign point_4_x[36] = 7'd6;
assign point_4_y[36] = 7'd50;
assign point_4_x[37] = 7'd5;
assign point_4_y[37] = 7'd47;
assign point_4_x[38] = 7'd6;
assign point_4_y[38] = 7'd43;
assign point_4_x[39] = 7'd6;
assign point_4_y[39] = 7'd40;
assign point_4_x[40] = 7'd8;
assign point_4_y[40] = 7'd36;
assign point_4_x[41] = 7'd9;
assign point_4_y[41] = 7'd33;
assign point_4_x[42] = 7'd12;
assign point_4_y[42] = 7'd29;
assign point_4_x[43] = 7'd15;
assign point_4_y[43] = 7'd25;
assign point_4_x[44] = 7'd18;
assign point_4_y[44] = 7'd22;
assign point_4_x[45] = 7'd22;
assign point_4_y[45] = 7'd18;
assign point_4_x[46] = 7'd26;
assign point_4_y[46] = 7'd15;
assign point_4_x[47] = 7'd30;
assign point_4_y[47] = 7'd13;
assign point_4_x[48] = 7'd35;
assign point_4_y[48] = 7'd10;
assign point_4_x[49] = 7'd40;
assign point_4_y[49] = 7'd8;
assign point_4_x[50] = 7'd45;
assign point_4_y[50] = 7'd6;
assign point_4_x[51] = 7'd50;
assign point_4_y[51] = 7'd5;
assign point_4_x[52] = 7'd54;
assign point_4_y[52] = 7'd4;
assign point_4_x[53] = 7'd59;
assign point_4_y[53] = 7'd4;
assign point_4_x[54] = 7'd64;
assign point_4_y[54] = 7'd4;
assign point_4_x[55] = 7'd68;
assign point_4_y[55] = 7'd4;
assign point_4_x[56] = 7'd71;
assign point_4_y[56] = 7'd5;
assign point_4_x[57] = 7'd74;
assign point_4_y[57] = 7'd6;
assign point_4_x[58] = 7'd77;
assign point_4_y[58] = 7'd7;
assign point_4_x[59] = 7'd79;
assign point_4_y[59] = 7'd8;
assign point_4_x[60] = 7'd80;
assign point_4_y[60] = 7'd10;
assign point_4_x[61] = 7'd81;
assign point_4_y[61] = 7'd11;
assign point_4_x[62] = 7'd81;
assign point_4_y[62] = 7'd13;
assign point_4_x[63] = 7'd81;
assign point_4_y[63] = 7'd15;
logic [types::LINE_BITS-1:0] point_5_x [64];
logic [types::LINE_BITS-1:0] point_5_y [64];
assign point_5_x[0] = 7'd80;
assign point_5_y[0] = 7'd59;
assign point_5_x[1] = 7'd75;
assign point_5_y[1] = 7'd60;
assign point_5_x[2] = 7'd70;
assign point_5_y[2] = 7'd61;
assign point_5_x[3] = 7'd66;
assign point_5_y[3] = 7'd62;
assign point_5_x[4] = 7'd61;
assign point_5_y[4] = 7'd62;
assign point_5_x[5] = 7'd56;
assign point_5_y[5] = 7'd63;
assign point_5_x[6] = 7'd51;
assign point_5_y[6] = 7'd63;
assign point_5_x[7] = 7'd46;
assign point_5_y[7] = 7'd62;
assign point_5_x[8] = 7'd42;
assign point_5_y[8] = 7'd62;
assign point_5_x[9] = 7'd37;
assign point_5_y[9] = 7'd61;
assign point_5_x[10] = 7'd33;
assign point_5_y[10] = 7'd59;
assign point_5_x[11] = 7'd29;
assign point_5_y[11] = 7'd58;
assign point_5_x[12] = 7'd25;
assign point_5_y[12] = 7'd57;
assign point_5_x[13] = 7'd21;
assign point_5_y[13] = 7'd55;
assign point_5_x[14] = 7'd18;
assign point_5_y[14] = 7'd53;
assign point_5_x[15] = 7'd15;
assign point_5_y[15] = 7'd51;
assign point_5_x[16] = 7'd13;
assign point_5_y[16] = 7'd49;
assign point_5_x[17] = 7'd10;
assign point_5_y[17] = 7'd47;
assign point_5_x[18] = 7'd8;
assign point_5_y[18] = 7'd44;
assign point_5_x[19] = 7'd7;
assign point_5_y[19] = 7'd42;
assign point_5_x[20] = 7'd6;
assign point_5_y[20] = 7'd40;
assign point_5_x[21] = 7'd5;
assign point_5_y[21] = 7'd38;
assign point_5_x[22] = 7'd4;
assign point_5_y[22] = 7'd35;
assign point_5_x[23] = 7'd3;
assign point_5_y[23] = 7'd33;
assign point_5_x[24] = 7'd3;
assign point_5_y[24] = 7'd31;
assign point_5_x[25] = 7'd3;
assign point_5_y[25] = 7'd29;
assign point_5_x[26] = 7'd4;
assign point_5_y[26] = 7'd27;
assign point_5_x[27] = 7'd4;
assign point_5_y[27] = 7'd25;
assign point_5_x[28] = 7'd5;
assign point_5_y[28] = 7'd23;
assign point_5_x[29] = 7'd6;
assign point_5_y[29] = 7'd21;
assign point_5_x[30] = 7'd7;
assign point_5_y[30] = 7'd20;
assign point_5_x[31] = 7'd8;
assign point_5_y[31] = 7'd18;
assign point_5_x[32] = 7'd9;
assign point_5_y[32] = 7'd16;
assign point_5_x[33] = 7'd11;
assign point_5_y[33] = 7'd15;
assign point_5_x[34] = 7'd13;
assign point_5_y[34] = 7'd14;
assign point_5_x[35] = 7'd14;
assign point_5_y[35] = 7'd13;
assign point_5_x[36] = 7'd16;
assign point_5_y[36] = 7'd12;
assign point_5_x[37] = 7'd18;
assign point_5_y[37] = 7'd11;
assign point_5_x[38] = 7'd20;
assign point_5_y[38] = 7'd10;
assign point_5_x[39] = 7'd22;
assign point_5_y[39] = 7'd9;
assign point_5_x[40] = 7'd23;
assign point_5_y[40] = 7'd9;
assign point_5_x[41] = 7'd25;
assign point_5_y[41] = 7'd9;
assign point_5_x[42] = 7'd27;
assign point_5_y[42] = 7'd8;
assign point_5_x[43] = 7'd29;
assign point_5_y[43] = 7'd8;
assign point_5_x[44] = 7'd30;
assign point_5_y[44] = 7'd8;
assign point_5_x[45] = 7'd32;
assign point_5_y[45] = 7'd9;
assign point_5_x[46] = 7'd33;
assign point_5_y[46] = 7'd9;
assign point_5_x[47] = 7'd34;
assign point_5_y[47] = 7'd9;
assign point_5_x[48] = 7'd35;
assign point_5_y[48] = 7'd10;
assign point_5_x[49] = 7'd35;
assign point_5_y[49] = 7'd11;
assign point_5_x[50] = 7'd36;
assign point_5_y[50] = 7'd11;
assign point_5_x[51] = 7'd36;
assign point_5_y[51] = 7'd12;
assign point_5_x[52] = 7'd36;
assign point_5_y[52] = 7'd13;
assign point_5_x[53] = 7'd36;
assign point_5_y[53] = 7'd14;
assign point_5_x[54] = 7'd35;
assign point_5_y[54] = 7'd15;
assign point_5_x[55] = 7'd34;
assign point_5_y[55] = 7'd15;
assign point_5_x[56] = 7'd33;
assign point_5_y[56] = 7'd16;
assign point_5_x[57] = 7'd32;
assign point_5_y[57] = 7'd16;
assign point_5_x[58] = 7'd31;
assign point_5_y[58] = 7'd17;
assign point_5_x[59] = 7'd29;
assign point_5_y[59] = 7'd17;
assign point_5_x[60] = 7'd28;
assign point_5_y[60] = 7'd17;
assign point_5_x[61] = 7'd26;
assign point_5_y[61] = 7'd17;
assign point_5_x[62] = 7'd25;
assign point_5_y[62] = 7'd17;
assign point_5_x[63] = 7'd23;
assign point_5_y[63] = 7'd17;
logic [types::LINE_BITS-1:0] point_6_x [64];
logic [types::LINE_BITS-1:0] point_6_y [64];
assign point_6_x[0] = 7'd22;
assign point_6_y[0] = 7'd59;
assign point_6_x[1] = 7'd23;
assign point_6_y[1] = 7'd57;
assign point_6_x[2] = 7'd25;
assign point_6_y[2] = 7'd56;
assign point_6_x[3] = 7'd28;
assign point_6_y[3] = 7'd55;
assign point_6_x[4] = 7'd31;
assign point_6_y[4] = 7'd54;
assign point_6_x[5] = 7'd34;
assign point_6_y[5] = 7'd53;
assign point_6_x[6] = 7'd38;
assign point_6_y[6] = 7'd53;
assign point_6_x[7] = 7'd41;
assign point_6_y[7] = 7'd53;
assign point_6_x[8] = 7'd45;
assign point_6_y[8] = 7'd54;
assign point_6_x[9] = 7'd49;
assign point_6_y[9] = 7'd54;
assign point_6_x[10] = 7'd52;
assign point_6_y[10] = 7'd55;
assign point_6_x[11] = 7'd55;
assign point_6_y[11] = 7'd57;
assign point_6_x[12] = 7'd58;
assign point_6_y[12] = 7'd58;
assign point_6_x[13] = 7'd61;
assign point_6_y[13] = 7'd60;
assign point_6_x[14] = 7'd63;
assign point_6_y[14] = 7'd61;
assign point_6_x[15] = 7'd65;
assign point_6_y[15] = 7'd63;
assign point_6_x[16] = 7'd66;
assign point_6_y[16] = 7'd65;
assign point_6_x[17] = 7'd67;
assign point_6_y[17] = 7'd67;
assign point_6_x[18] = 7'd67;
assign point_6_y[18] = 7'd68;
assign point_6_x[19] = 7'd67;
assign point_6_y[19] = 7'd70;
assign point_6_x[20] = 7'd67;
assign point_6_y[20] = 7'd71;
assign point_6_x[21] = 7'd66;
assign point_6_y[21] = 7'd72;
assign point_6_x[22] = 7'd65;
assign point_6_y[22] = 7'd72;
assign point_6_x[23] = 7'd63;
assign point_6_y[23] = 7'd73;
assign point_6_x[24] = 7'd62;
assign point_6_y[24] = 7'd72;
assign point_6_x[25] = 7'd60;
assign point_6_y[25] = 7'd72;
assign point_6_x[26] = 7'd58;
assign point_6_y[26] = 7'd71;
assign point_6_x[27] = 7'd57;
assign point_6_y[27] = 7'd70;
assign point_6_x[28] = 7'd55;
assign point_6_y[28] = 7'd68;
assign point_6_x[29] = 7'd53;
assign point_6_y[29] = 7'd66;
assign point_6_x[30] = 7'd52;
assign point_6_y[30] = 7'd64;
assign point_6_x[31] = 7'd51;
assign point_6_y[31] = 7'd61;
assign point_6_x[32] = 7'd50;
assign point_6_y[32] = 7'd58;
assign point_6_x[33] = 7'd50;
assign point_6_y[33] = 7'd56;
assign point_6_x[34] = 7'd50;
assign point_6_y[34] = 7'd52;
assign point_6_x[35] = 7'd51;
assign point_6_y[35] = 7'd49;
assign point_6_x[36] = 7'd52;
assign point_6_y[36] = 7'd46;
assign point_6_x[37] = 7'd54;
assign point_6_y[37] = 7'd43;
assign point_6_x[38] = 7'd56;
assign point_6_y[38] = 7'd40;
assign point_6_x[39] = 7'd58;
assign point_6_y[39] = 7'd37;
assign point_6_x[40] = 7'd61;
assign point_6_y[40] = 7'd34;
assign point_6_x[41] = 7'd64;
assign point_6_y[41] = 7'd32;
assign point_6_x[42] = 7'd67;
assign point_6_y[42] = 7'd30;
assign point_6_x[43] = 7'd71;
assign point_6_y[43] = 7'd28;
assign point_6_x[44] = 7'd74;
assign point_6_y[44] = 7'd27;
assign point_6_x[45] = 7'd78;
assign point_6_y[45] = 7'd26;
assign point_6_x[46] = 7'd82;
assign point_6_y[46] = 7'd26;
assign point_6_x[47] = 7'd85;
assign point_6_y[47] = 7'd26;
assign point_6_x[48] = 7'd88;
assign point_6_y[48] = 7'd26;
assign point_6_x[49] = 7'd91;
assign point_6_y[49] = 7'd27;
assign point_6_x[50] = 7'd94;
assign point_6_y[50] = 7'd28;
assign point_6_x[51] = 7'd96;
assign point_6_y[51] = 7'd29;
assign point_6_x[52] = 7'd98;
assign point_6_y[52] = 7'd31;
assign point_6_x[53] = 7'd100;
assign point_6_y[53] = 7'd33;
assign point_6_x[54] = 7'd100;
assign point_6_y[54] = 7'd35;
assign point_6_x[55] = 7'd101;
assign point_6_y[55] = 7'd38;
assign point_6_x[56] = 7'd100;
assign point_6_y[56] = 7'd40;
assign point_6_x[57] = 7'd100;
assign point_6_y[57] = 7'd43;
assign point_6_x[58] = 7'd98;
assign point_6_y[58] = 7'd46;
assign point_6_x[59] = 7'd96;
assign point_6_y[59] = 7'd48;
assign point_6_x[60] = 7'd94;
assign point_6_y[60] = 7'd50;
assign point_6_x[61] = 7'd91;
assign point_6_y[61] = 7'd53;
assign point_6_x[62] = 7'd87;
assign point_6_y[62] = 7'd55;
assign point_6_x[63] = 7'd84;
assign point_6_y[63] = 7'd57;
logic [types::LINE_BITS-1:0] point_7_x [64];
logic [types::LINE_BITS-1:0] point_7_y [64];
assign point_7_x[0] = 7'd80;
assign point_7_y[0] = 7'd59;
assign point_7_x[1] = 7'd81;
assign point_7_y[1] = 7'd59;
assign point_7_x[2] = 7'd82;
assign point_7_y[2] = 7'd60;
assign point_7_x[3] = 7'd83;
assign point_7_y[3] = 7'd61;
assign point_7_x[4] = 7'd84;
assign point_7_y[4] = 7'd61;
assign point_7_x[5] = 7'd84;
assign point_7_y[5] = 7'd62;
assign point_7_x[6] = 7'd84;
assign point_7_y[6] = 7'd63;
assign point_7_x[7] = 7'd84;
assign point_7_y[7] = 7'd64;
assign point_7_x[8] = 7'd83;
assign point_7_y[8] = 7'd65;
assign point_7_x[9] = 7'd82;
assign point_7_y[9] = 7'd66;
assign point_7_x[10] = 7'd81;
assign point_7_y[10] = 7'd66;
assign point_7_x[11] = 7'd79;
assign point_7_y[11] = 7'd67;
assign point_7_x[12] = 7'd77;
assign point_7_y[12] = 7'd67;
assign point_7_x[13] = 7'd74;
assign point_7_y[13] = 7'd67;
assign point_7_x[14] = 7'd72;
assign point_7_y[14] = 7'd67;
assign point_7_x[15] = 7'd69;
assign point_7_y[15] = 7'd66;
assign point_7_x[16] = 7'd66;
assign point_7_y[16] = 7'd65;
assign point_7_x[17] = 7'd63;
assign point_7_y[17] = 7'd64;
assign point_7_x[18] = 7'd60;
assign point_7_y[18] = 7'd62;
assign point_7_x[19] = 7'd57;
assign point_7_y[19] = 7'd60;
assign point_7_x[20] = 7'd55;
assign point_7_y[20] = 7'd57;
assign point_7_x[21] = 7'd52;
assign point_7_y[21] = 7'd55;
assign point_7_x[22] = 7'd50;
assign point_7_y[22] = 7'd52;
assign point_7_x[23] = 7'd48;
assign point_7_y[23] = 7'd48;
assign point_7_x[24] = 7'd46;
assign point_7_y[24] = 7'd45;
assign point_7_x[25] = 7'd45;
assign point_7_y[25] = 7'd41;
assign point_7_x[26] = 7'd44;
assign point_7_y[26] = 7'd38;
assign point_7_x[27] = 7'd44;
assign point_7_y[27] = 7'd34;
assign point_7_x[28] = 7'd44;
assign point_7_y[28] = 7'd30;
assign point_7_x[29] = 7'd45;
assign point_7_y[29] = 7'd26;
assign point_7_x[30] = 7'd46;
assign point_7_y[30] = 7'd23;
assign point_7_x[31] = 7'd48;
assign point_7_y[31] = 7'd20;
assign point_7_x[32] = 7'd51;
assign point_7_y[32] = 7'd16;
assign point_7_x[33] = 7'd53;
assign point_7_y[33] = 7'd14;
assign point_7_x[34] = 7'd56;
assign point_7_y[34] = 7'd11;
assign point_7_x[35] = 7'd59;
assign point_7_y[35] = 7'd9;
assign point_7_x[36] = 7'd63;
assign point_7_y[36] = 7'd8;
assign point_7_x[37] = 7'd66;
assign point_7_y[37] = 7'd7;
assign point_7_x[38] = 7'd70;
assign point_7_y[38] = 7'd6;
assign point_7_x[39] = 7'd73;
assign point_7_y[39] = 7'd6;
assign point_7_x[40] = 7'd77;
assign point_7_y[40] = 7'd7;
assign point_7_x[41] = 7'd80;
assign point_7_y[41] = 7'd8;
assign point_7_x[42] = 7'd82;
assign point_7_y[42] = 7'd9;
assign point_7_x[43] = 7'd85;
assign point_7_y[43] = 7'd11;
assign point_7_x[44] = 7'd87;
assign point_7_y[44] = 7'd14;
assign point_7_x[45] = 7'd88;
assign point_7_y[45] = 7'd16;
assign point_7_x[46] = 7'd89;
assign point_7_y[46] = 7'd19;
assign point_7_x[47] = 7'd89;
assign point_7_y[47] = 7'd23;
assign point_7_x[48] = 7'd88;
assign point_7_y[48] = 7'd26;
assign point_7_x[49] = 7'd87;
assign point_7_y[49] = 7'd30;
assign point_7_x[50] = 7'd85;
assign point_7_y[50] = 7'd33;
assign point_7_x[51] = 7'd83;
assign point_7_y[51] = 7'd37;
assign point_7_x[52] = 7'd80;
assign point_7_y[52] = 7'd40;
assign point_7_x[53] = 7'd76;
assign point_7_y[53] = 7'd43;
assign point_7_x[54] = 7'd72;
assign point_7_y[54] = 7'd46;
assign point_7_x[55] = 7'd67;
assign point_7_y[55] = 7'd49;
assign point_7_x[56] = 7'd63;
assign point_7_y[56] = 7'd52;
assign point_7_x[57] = 7'd57;
assign point_7_y[57] = 7'd54;
assign point_7_x[58] = 7'd52;
assign point_7_y[58] = 7'd56;
assign point_7_x[59] = 7'd47;
assign point_7_y[59] = 7'd57;
assign point_7_x[60] = 7'd41;
assign point_7_y[60] = 7'd58;
assign point_7_x[61] = 7'd36;
assign point_7_y[61] = 7'd59;
assign point_7_x[62] = 7'd31;
assign point_7_y[62] = 7'd59;
assign point_7_x[63] = 7'd26;
assign point_7_y[63] = 7'd59;
logic [types::THRESH_BITS-1:0] threshold_0 [64];
assign threshold_0[0] = 8'd58;
assign threshold_0[1] = 8'd58;
assign threshold_0[2] = 8'd57;
assign threshold_0[3] = 8'd55;
assign threshold_0[4] = 8'd53;
assign threshold_0[5] = 8'd51;
assign threshold_0[6] = 8'd47;
assign threshold_0[7] = 8'd44;
assign threshold_0[8] = 8'd40;
assign threshold_0[9] = 8'd35;
assign threshold_0[10] = 8'd31;
assign threshold_0[11] = 8'd26;
assign threshold_0[12] = 8'd21;
assign threshold_0[13] = 8'd15;
assign threshold_0[14] = 8'd11;
assign threshold_0[15] = 8'd5;
assign threshold_0[16] = 8'd0;
assign threshold_0[17] = 8'd5;
assign threshold_0[18] = 8'd9;
assign threshold_0[19] = 8'd14;
assign threshold_0[20] = 8'd18;
assign threshold_0[21] = 8'd22;
assign threshold_0[22] = 8'd25;
assign threshold_0[23] = 8'd29;
assign threshold_0[24] = 8'd31;
assign threshold_0[25] = 8'd34;
assign threshold_0[26] = 8'd36;
assign threshold_0[27] = 8'd38;
assign threshold_0[28] = 8'd40;
assign threshold_0[29] = 8'd41;
assign threshold_0[30] = 8'd41;
assign threshold_0[31] = 8'd41;
assign threshold_0[32] = 8'd42;
assign threshold_0[33] = 8'd42;
assign threshold_0[34] = 8'd41;
assign threshold_0[35] = 8'd41;
assign threshold_0[36] = 8'd40;
assign threshold_0[37] = 8'd38;
assign threshold_0[38] = 8'd37;
assign threshold_0[39] = 8'd34;
assign threshold_0[40] = 8'd31;
assign threshold_0[41] = 8'd29;
assign threshold_0[42] = 8'd26;
assign threshold_0[43] = 8'd22;
assign threshold_0[44] = 8'd18;
assign threshold_0[45] = 8'd14;
assign threshold_0[46] = 8'd10;
assign threshold_0[47] = 8'd5;
assign threshold_0[48] = 8'd0;
assign threshold_0[49] = 8'd5;
assign threshold_0[50] = 8'd10;
assign threshold_0[51] = 8'd15;
assign threshold_0[52] = 8'd20;
assign threshold_0[53] = 8'd26;
assign threshold_0[54] = 8'd30;
assign threshold_0[55] = 8'd36;
assign threshold_0[56] = 8'd39;
assign threshold_0[57] = 8'd44;
assign threshold_0[58] = 8'd47;
assign threshold_0[59] = 8'd50;
assign threshold_0[60] = 8'd54;
assign threshold_0[61] = 8'd55;
assign threshold_0[62] = 8'd56;
assign threshold_0[63] = 8'd58;
logic [types::THRESH_BITS-1:0] threshold_1 [64];
assign threshold_1[0] = 8'd0;
assign threshold_1[1] = 8'd6;
assign threshold_1[2] = 8'd11;
assign threshold_1[3] = 8'd17;
assign threshold_1[4] = 8'd23;
assign threshold_1[5] = 8'd28;
assign threshold_1[6] = 8'd33;
assign threshold_1[7] = 8'd37;
assign threshold_1[8] = 8'd41;
assign threshold_1[9] = 8'd45;
assign threshold_1[10] = 8'd49;
assign threshold_1[11] = 8'd51;
assign threshold_1[12] = 8'd53;
assign threshold_1[13] = 8'd54;
assign threshold_1[14] = 8'd56;
assign threshold_1[15] = 8'd56;
assign threshold_1[16] = 8'd55;
assign threshold_1[17] = 8'd56;
assign threshold_1[18] = 8'd54;
assign threshold_1[19] = 8'd53;
assign threshold_1[20] = 8'd52;
assign threshold_1[21] = 8'd50;
assign threshold_1[22] = 8'd49;
assign threshold_1[23] = 8'd47;
assign threshold_1[24] = 8'd45;
assign threshold_1[25] = 8'd43;
assign threshold_1[26] = 8'd41;
assign threshold_1[27] = 8'd41;
assign threshold_1[28] = 8'd41;
assign threshold_1[29] = 8'd39;
assign threshold_1[30] = 8'd40;
assign threshold_1[31] = 8'd40;
assign threshold_1[32] = 8'd41;
assign threshold_1[33] = 8'd42;
assign threshold_1[34] = 8'd43;
assign threshold_1[35] = 8'd45;
assign threshold_1[36] = 8'd46;
assign threshold_1[37] = 8'd49;
assign threshold_1[38] = 8'd50;
assign threshold_1[39] = 8'd52;
assign threshold_1[40] = 8'd53;
assign threshold_1[41] = 8'd55;
assign threshold_1[42] = 8'd55;
assign threshold_1[43] = 8'd56;
assign threshold_1[44] = 8'd56;
assign threshold_1[45] = 8'd57;
assign threshold_1[46] = 8'd57;
assign threshold_1[47] = 8'd57;
assign threshold_1[48] = 8'd55;
assign threshold_1[49] = 8'd54;
assign threshold_1[50] = 8'd54;
assign threshold_1[51] = 8'd52;
assign threshold_1[52] = 8'd52;
assign threshold_1[53] = 8'd50;
assign threshold_1[54] = 8'd48;
assign threshold_1[55] = 8'd47;
assign threshold_1[56] = 8'd45;
assign threshold_1[57] = 8'd45;
assign threshold_1[58] = 8'd44;
assign threshold_1[59] = 8'd43;
assign threshold_1[60] = 8'd42;
assign threshold_1[61] = 8'd43;
assign threshold_1[62] = 8'd42;
assign threshold_1[63] = 8'd42;
logic [types::THRESH_BITS-1:0] threshold_2 [64];
assign threshold_2[0] = 8'd58;
assign threshold_2[1] = 8'd58;
assign threshold_2[2] = 8'd56;
assign threshold_2[3] = 8'd55;
assign threshold_2[4] = 8'd53;
assign threshold_2[5] = 8'd51;
assign threshold_2[6] = 8'd47;
assign threshold_2[7] = 8'd43;
assign threshold_2[8] = 8'd40;
assign threshold_2[9] = 8'd35;
assign threshold_2[10] = 8'd31;
assign threshold_2[11] = 8'd26;
assign threshold_2[12] = 8'd21;
assign threshold_2[13] = 8'd15;
assign threshold_2[14] = 8'd10;
assign threshold_2[15] = 8'd5;
assign threshold_2[16] = 8'd0;
assign threshold_2[17] = 8'd5;
assign threshold_2[18] = 8'd11;
assign threshold_2[19] = 8'd14;
assign threshold_2[20] = 8'd18;
assign threshold_2[21] = 8'd22;
assign threshold_2[22] = 8'd26;
assign threshold_2[23] = 8'd29;
assign threshold_2[24] = 8'd32;
assign threshold_2[25] = 8'd35;
assign threshold_2[26] = 8'd36;
assign threshold_2[27] = 8'd38;
assign threshold_2[28] = 8'd39;
assign threshold_2[29] = 8'd41;
assign threshold_2[30] = 8'd41;
assign threshold_2[31] = 8'd42;
assign threshold_2[32] = 8'd42;
assign threshold_2[33] = 8'd42;
assign threshold_2[34] = 8'd41;
assign threshold_2[35] = 8'd40;
assign threshold_2[36] = 8'd39;
assign threshold_2[37] = 8'd38;
assign threshold_2[38] = 8'd36;
assign threshold_2[39] = 8'd35;
assign threshold_2[40] = 8'd31;
assign threshold_2[41] = 8'd29;
assign threshold_2[42] = 8'd26;
assign threshold_2[43] = 8'd22;
assign threshold_2[44] = 8'd18;
assign threshold_2[45] = 8'd13;
assign threshold_2[46] = 8'd9;
assign threshold_2[47] = 8'd6;
assign threshold_2[48] = 8'd0;
assign threshold_2[49] = 8'd6;
assign threshold_2[50] = 8'd10;
assign threshold_2[51] = 8'd16;
assign threshold_2[52] = 8'd20;
assign threshold_2[53] = 8'd25;
assign threshold_2[54] = 8'd31;
assign threshold_2[55] = 8'd36;
assign threshold_2[56] = 8'd40;
assign threshold_2[57] = 8'd43;
assign threshold_2[58] = 8'd47;
assign threshold_2[59] = 8'd51;
assign threshold_2[60] = 8'd52;
assign threshold_2[61] = 8'd55;
assign threshold_2[62] = 8'd56;
assign threshold_2[63] = 8'd58;
logic [types::THRESH_BITS-1:0] threshold_3 [64];
assign threshold_3[0] = 8'd0;
assign threshold_3[1] = 8'd6;
assign threshold_3[2] = 8'd12;
assign threshold_3[3] = 8'd17;
assign threshold_3[4] = 8'd23;
assign threshold_3[5] = 8'd28;
assign threshold_3[6] = 8'd33;
assign threshold_3[7] = 8'd38;
assign threshold_3[8] = 8'd41;
assign threshold_3[9] = 8'd45;
assign threshold_3[10] = 8'd49;
assign threshold_3[11] = 8'd51;
assign threshold_3[12] = 8'd53;
assign threshold_3[13] = 8'd54;
assign threshold_3[14] = 8'd56;
assign threshold_3[15] = 8'd56;
assign threshold_3[16] = 8'd55;
assign threshold_3[17] = 8'd56;
assign threshold_3[18] = 8'd55;
assign threshold_3[19] = 8'd53;
assign threshold_3[20] = 8'd52;
assign threshold_3[21] = 8'd50;
assign threshold_3[22] = 8'd49;
assign threshold_3[23] = 8'd47;
assign threshold_3[24] = 8'd45;
assign threshold_3[25] = 8'd44;
assign threshold_3[26] = 8'd41;
assign threshold_3[27] = 8'd41;
assign threshold_3[28] = 8'd40;
assign threshold_3[29] = 8'd39;
assign threshold_3[30] = 8'd39;
assign threshold_3[31] = 8'd40;
assign threshold_3[32] = 8'd42;
assign threshold_3[33] = 8'd42;
assign threshold_3[34] = 8'd43;
assign threshold_3[35] = 8'd45;
assign threshold_3[36] = 8'd47;
assign threshold_3[37] = 8'd48;
assign threshold_3[38] = 8'd50;
assign threshold_3[39] = 8'd51;
assign threshold_3[40] = 8'd54;
assign threshold_3[41] = 8'd55;
assign threshold_3[42] = 8'd55;
assign threshold_3[43] = 8'd56;
assign threshold_3[44] = 8'd57;
assign threshold_3[45] = 8'd56;
assign threshold_3[46] = 8'd57;
assign threshold_3[47] = 8'd57;
assign threshold_3[48] = 8'd55;
assign threshold_3[49] = 8'd55;
assign threshold_3[50] = 8'd54;
assign threshold_3[51] = 8'd53;
assign threshold_3[52] = 8'd52;
assign threshold_3[53] = 8'd49;
assign threshold_3[54] = 8'd48;
assign threshold_3[55] = 8'd47;
assign threshold_3[56] = 8'd47;
assign threshold_3[57] = 8'd45;
assign threshold_3[58] = 8'd44;
assign threshold_3[59] = 8'd44;
assign threshold_3[60] = 8'd43;
assign threshold_3[61] = 8'd43;
assign threshold_3[62] = 8'd42;
assign threshold_3[63] = 8'd42;
logic [types::THRESH_BITS-1:0] threshold_4 [64];
assign threshold_4[0] = 8'd42;
assign threshold_4[1] = 8'd42;
assign threshold_4[2] = 8'd42;
assign threshold_4[3] = 8'd43;
assign threshold_4[4] = 8'd42;
assign threshold_4[5] = 8'd42;
assign threshold_4[6] = 8'd42;
assign threshold_4[7] = 8'd42;
assign threshold_4[8] = 8'd42;
assign threshold_4[9] = 8'd43;
assign threshold_4[10] = 8'd42;
assign threshold_4[11] = 8'd43;
assign threshold_4[12] = 8'd44;
assign threshold_4[13] = 8'd44;
assign threshold_4[14] = 8'd45;
assign threshold_4[15] = 8'd44;
assign threshold_4[16] = 8'd45;
assign threshold_4[17] = 8'd46;
assign threshold_4[18] = 8'd45;
assign threshold_4[19] = 8'd46;
assign threshold_4[20] = 8'd45;
assign threshold_4[21] = 8'd46;
assign threshold_4[22] = 8'd46;
assign threshold_4[23] = 8'd45;
assign threshold_4[24] = 8'd46;
assign threshold_4[25] = 8'd45;
assign threshold_4[26] = 8'd45;
assign threshold_4[27] = 8'd45;
assign threshold_4[28] = 8'd45;
assign threshold_4[29] = 8'd44;
assign threshold_4[30] = 8'd44;
assign threshold_4[31] = 8'd42;
assign threshold_4[32] = 8'd41;
assign threshold_4[33] = 8'd40;
assign threshold_4[34] = 8'd39;
assign threshold_4[35] = 8'd39;
assign threshold_4[36] = 8'd36;
assign threshold_4[37] = 8'd37;
assign threshold_4[38] = 8'd36;
assign threshold_4[39] = 8'd36;
assign threshold_4[40] = 8'd36;
assign threshold_4[41] = 8'd36;
assign threshold_4[42] = 8'd38;
assign threshold_4[43] = 8'd39;
assign threshold_4[44] = 8'd39;
assign threshold_4[45] = 8'd42;
assign threshold_4[46] = 8'd43;
assign threshold_4[47] = 8'd43;
assign threshold_4[48] = 8'd45;
assign threshold_4[49] = 8'd45;
assign threshold_4[50] = 8'd46;
assign threshold_4[51] = 8'd46;
assign threshold_4[52] = 8'd45;
assign threshold_4[53] = 8'd44;
assign threshold_4[54] = 8'd43;
assign threshold_4[55] = 8'd40;
assign threshold_4[56] = 8'd38;
assign threshold_4[57] = 8'd34;
assign threshold_4[58] = 8'd30;
assign threshold_4[59] = 8'd27;
assign threshold_4[60] = 8'd21;
assign threshold_4[61] = 8'd17;
assign threshold_4[62] = 8'd11;
assign threshold_4[63] = 8'd6;
logic [types::THRESH_BITS-1:0] threshold_5 [64];
assign threshold_5[0] = 8'd42;
assign threshold_5[1] = 8'd42;
assign threshold_5[2] = 8'd42;
assign threshold_5[3] = 8'd43;
assign threshold_5[4] = 8'd42;
assign threshold_5[5] = 8'd42;
assign threshold_5[6] = 8'd43;
assign threshold_5[7] = 8'd42;
assign threshold_5[8] = 8'd43;
assign threshold_5[9] = 8'd43;
assign threshold_5[10] = 8'd42;
assign threshold_5[11] = 8'd43;
assign threshold_5[12] = 8'd44;
assign threshold_5[13] = 8'd44;
assign threshold_5[14] = 8'd44;
assign threshold_5[15] = 8'd44;
assign threshold_5[16] = 8'd45;
assign threshold_5[17] = 8'd46;
assign threshold_5[18] = 8'd45;
assign threshold_5[19] = 8'd46;
assign threshold_5[20] = 8'd46;
assign threshold_5[21] = 8'd46;
assign threshold_5[22] = 8'd45;
assign threshold_5[23] = 8'd47;
assign threshold_5[24] = 8'd46;
assign threshold_5[25] = 8'd46;
assign threshold_5[26] = 8'd45;
assign threshold_5[27] = 8'd45;
assign threshold_5[28] = 8'd44;
assign threshold_5[29] = 8'd44;
assign threshold_5[30] = 8'd43;
assign threshold_5[31] = 8'd42;
assign threshold_5[32] = 8'd42;
assign threshold_5[33] = 8'd40;
assign threshold_5[34] = 8'd39;
assign threshold_5[35] = 8'd38;
assign threshold_5[36] = 8'd37;
assign threshold_5[37] = 8'd36;
assign threshold_5[38] = 8'd35;
assign threshold_5[39] = 8'd36;
assign threshold_5[40] = 8'd36;
assign threshold_5[41] = 8'd36;
assign threshold_5[42] = 8'd38;
assign threshold_5[43] = 8'd39;
assign threshold_5[44] = 8'd40;
assign threshold_5[45] = 8'd41;
assign threshold_5[46] = 8'd42;
assign threshold_5[47] = 8'd44;
assign threshold_5[48] = 8'd45;
assign threshold_5[49] = 8'd45;
assign threshold_5[50] = 8'd46;
assign threshold_5[51] = 8'd46;
assign threshold_5[52] = 8'd45;
assign threshold_5[53] = 8'd45;
assign threshold_5[54] = 8'd42;
assign threshold_5[55] = 8'd40;
assign threshold_5[56] = 8'd37;
assign threshold_5[57] = 8'd35;
assign threshold_5[58] = 8'd30;
assign threshold_5[59] = 8'd26;
assign threshold_5[60] = 8'd22;
assign threshold_5[61] = 8'd17;
assign threshold_5[62] = 8'd11;
assign threshold_5[63] = 8'd6;
logic [types::THRESH_BITS-1:0] threshold_6 [64];
assign threshold_6[0] = 8'd42;
assign threshold_6[1] = 8'd42;
assign threshold_6[2] = 8'd42;
assign threshold_6[3] = 8'd43;
assign threshold_6[4] = 8'd42;
assign threshold_6[5] = 8'd42;
assign threshold_6[6] = 8'd43;
assign threshold_6[7] = 8'd42;
assign threshold_6[8] = 8'd43;
assign threshold_6[9] = 8'd43;
assign threshold_6[10] = 8'd42;
assign threshold_6[11] = 8'd43;
assign threshold_6[12] = 8'd44;
assign threshold_6[13] = 8'd44;
assign threshold_6[14] = 8'd44;
assign threshold_6[15] = 8'd44;
assign threshold_6[16] = 8'd45;
assign threshold_6[17] = 8'd46;
assign threshold_6[18] = 8'd45;
assign threshold_6[19] = 8'd46;
assign threshold_6[20] = 8'd46;
assign threshold_6[21] = 8'd46;
assign threshold_6[22] = 8'd45;
assign threshold_6[23] = 8'd47;
assign threshold_6[24] = 8'd46;
assign threshold_6[25] = 8'd46;
assign threshold_6[26] = 8'd45;
assign threshold_6[27] = 8'd45;
assign threshold_6[28] = 8'd44;
assign threshold_6[29] = 8'd44;
assign threshold_6[30] = 8'd43;
assign threshold_6[31] = 8'd42;
assign threshold_6[32] = 8'd42;
assign threshold_6[33] = 8'd40;
assign threshold_6[34] = 8'd39;
assign threshold_6[35] = 8'd38;
assign threshold_6[36] = 8'd37;
assign threshold_6[37] = 8'd36;
assign threshold_6[38] = 8'd35;
assign threshold_6[39] = 8'd36;
assign threshold_6[40] = 8'd36;
assign threshold_6[41] = 8'd36;
assign threshold_6[42] = 8'd38;
assign threshold_6[43] = 8'd39;
assign threshold_6[44] = 8'd40;
assign threshold_6[45] = 8'd41;
assign threshold_6[46] = 8'd42;
assign threshold_6[47] = 8'd44;
assign threshold_6[48] = 8'd45;
assign threshold_6[49] = 8'd45;
assign threshold_6[50] = 8'd46;
assign threshold_6[51] = 8'd46;
assign threshold_6[52] = 8'd45;
assign threshold_6[53] = 8'd45;
assign threshold_6[54] = 8'd42;
assign threshold_6[55] = 8'd40;
assign threshold_6[56] = 8'd37;
assign threshold_6[57] = 8'd35;
assign threshold_6[58] = 8'd30;
assign threshold_6[59] = 8'd26;
assign threshold_6[60] = 8'd22;
assign threshold_6[61] = 8'd17;
assign threshold_6[62] = 8'd11;
assign threshold_6[63] = 8'd6;
logic [types::THRESH_BITS-1:0] threshold_7 [64];
assign threshold_7[0] = 8'd42;
assign threshold_7[1] = 8'd42;
assign threshold_7[2] = 8'd42;
assign threshold_7[3] = 8'd43;
assign threshold_7[4] = 8'd42;
assign threshold_7[5] = 8'd42;
assign threshold_7[6] = 8'd42;
assign threshold_7[7] = 8'd42;
assign threshold_7[8] = 8'd42;
assign threshold_7[9] = 8'd43;
assign threshold_7[10] = 8'd42;
assign threshold_7[11] = 8'd43;
assign threshold_7[12] = 8'd44;
assign threshold_7[13] = 8'd44;
assign threshold_7[14] = 8'd45;
assign threshold_7[15] = 8'd44;
assign threshold_7[16] = 8'd45;
assign threshold_7[17] = 8'd46;
assign threshold_7[18] = 8'd45;
assign threshold_7[19] = 8'd46;
assign threshold_7[20] = 8'd45;
assign threshold_7[21] = 8'd46;
assign threshold_7[22] = 8'd46;
assign threshold_7[23] = 8'd45;
assign threshold_7[24] = 8'd46;
assign threshold_7[25] = 8'd45;
assign threshold_7[26] = 8'd45;
assign threshold_7[27] = 8'd45;
assign threshold_7[28] = 8'd45;
assign threshold_7[29] = 8'd44;
assign threshold_7[30] = 8'd44;
assign threshold_7[31] = 8'd42;
assign threshold_7[32] = 8'd41;
assign threshold_7[33] = 8'd40;
assign threshold_7[34] = 8'd39;
assign threshold_7[35] = 8'd39;
assign threshold_7[36] = 8'd36;
assign threshold_7[37] = 8'd37;
assign threshold_7[38] = 8'd36;
assign threshold_7[39] = 8'd36;
assign threshold_7[40] = 8'd36;
assign threshold_7[41] = 8'd36;
assign threshold_7[42] = 8'd38;
assign threshold_7[43] = 8'd39;
assign threshold_7[44] = 8'd39;
assign threshold_7[45] = 8'd42;
assign threshold_7[46] = 8'd43;
assign threshold_7[47] = 8'd43;
assign threshold_7[48] = 8'd45;
assign threshold_7[49] = 8'd45;
assign threshold_7[50] = 8'd46;
assign threshold_7[51] = 8'd46;
assign threshold_7[52] = 8'd45;
assign threshold_7[53] = 8'd44;
assign threshold_7[54] = 8'd43;
assign threshold_7[55] = 8'd40;
assign threshold_7[56] = 8'd38;
assign threshold_7[57] = 8'd34;
assign threshold_7[58] = 8'd30;
assign threshold_7[59] = 8'd27;
assign threshold_7[60] = 8'd21;
assign threshold_7[61] = 8'd17;
assign threshold_7[62] = 8'd11;
assign threshold_7[63] = 8'd6;
logic [types::THRESH_BITS-1:0] threshold_8 [64];
assign threshold_8[0] = 8'd58;
assign threshold_8[1] = 8'd58;
assign threshold_8[2] = 8'd56;
assign threshold_8[3] = 8'd55;
assign threshold_8[4] = 8'd53;
assign threshold_8[5] = 8'd51;
assign threshold_8[6] = 8'd47;
assign threshold_8[7] = 8'd43;
assign threshold_8[8] = 8'd40;
assign threshold_8[9] = 8'd35;
assign threshold_8[10] = 8'd31;
assign threshold_8[11] = 8'd26;
assign threshold_8[12] = 8'd21;
assign threshold_8[13] = 8'd15;
assign threshold_8[14] = 8'd10;
assign threshold_8[15] = 8'd5;
assign threshold_8[16] = 8'd0;
assign threshold_8[17] = 8'd5;
assign threshold_8[18] = 8'd11;
assign threshold_8[19] = 8'd14;
assign threshold_8[20] = 8'd18;
assign threshold_8[21] = 8'd22;
assign threshold_8[22] = 8'd26;
assign threshold_8[23] = 8'd29;
assign threshold_8[24] = 8'd32;
assign threshold_8[25] = 8'd35;
assign threshold_8[26] = 8'd36;
assign threshold_8[27] = 8'd38;
assign threshold_8[28] = 8'd39;
assign threshold_8[29] = 8'd41;
assign threshold_8[30] = 8'd41;
assign threshold_8[31] = 8'd42;
assign threshold_8[32] = 8'd42;
assign threshold_8[33] = 8'd42;
assign threshold_8[34] = 8'd41;
assign threshold_8[35] = 8'd40;
assign threshold_8[36] = 8'd39;
assign threshold_8[37] = 8'd38;
assign threshold_8[38] = 8'd36;
assign threshold_8[39] = 8'd35;
assign threshold_8[40] = 8'd31;
assign threshold_8[41] = 8'd29;
assign threshold_8[42] = 8'd26;
assign threshold_8[43] = 8'd22;
assign threshold_8[44] = 8'd18;
assign threshold_8[45] = 8'd13;
assign threshold_8[46] = 8'd9;
assign threshold_8[47] = 8'd6;
assign threshold_8[48] = 8'd0;
assign threshold_8[49] = 8'd6;
assign threshold_8[50] = 8'd10;
assign threshold_8[51] = 8'd16;
assign threshold_8[52] = 8'd20;
assign threshold_8[53] = 8'd25;
assign threshold_8[54] = 8'd31;
assign threshold_8[55] = 8'd36;
assign threshold_8[56] = 8'd40;
assign threshold_8[57] = 8'd43;
assign threshold_8[58] = 8'd47;
assign threshold_8[59] = 8'd51;
assign threshold_8[60] = 8'd52;
assign threshold_8[61] = 8'd55;
assign threshold_8[62] = 8'd56;
assign threshold_8[63] = 8'd58;
logic [types::THRESH_BITS-1:0] threshold_9 [64];
assign threshold_9[0] = 8'd0;
assign threshold_9[1] = 8'd6;
assign threshold_9[2] = 8'd12;
assign threshold_9[3] = 8'd17;
assign threshold_9[4] = 8'd23;
assign threshold_9[5] = 8'd28;
assign threshold_9[6] = 8'd33;
assign threshold_9[7] = 8'd38;
assign threshold_9[8] = 8'd41;
assign threshold_9[9] = 8'd45;
assign threshold_9[10] = 8'd49;
assign threshold_9[11] = 8'd51;
assign threshold_9[12] = 8'd53;
assign threshold_9[13] = 8'd54;
assign threshold_9[14] = 8'd56;
assign threshold_9[15] = 8'd56;
assign threshold_9[16] = 8'd55;
assign threshold_9[17] = 8'd56;
assign threshold_9[18] = 8'd55;
assign threshold_9[19] = 8'd53;
assign threshold_9[20] = 8'd52;
assign threshold_9[21] = 8'd50;
assign threshold_9[22] = 8'd49;
assign threshold_9[23] = 8'd47;
assign threshold_9[24] = 8'd45;
assign threshold_9[25] = 8'd44;
assign threshold_9[26] = 8'd41;
assign threshold_9[27] = 8'd41;
assign threshold_9[28] = 8'd40;
assign threshold_9[29] = 8'd39;
assign threshold_9[30] = 8'd39;
assign threshold_9[31] = 8'd40;
assign threshold_9[32] = 8'd42;
assign threshold_9[33] = 8'd42;
assign threshold_9[34] = 8'd43;
assign threshold_9[35] = 8'd45;
assign threshold_9[36] = 8'd47;
assign threshold_9[37] = 8'd48;
assign threshold_9[38] = 8'd50;
assign threshold_9[39] = 8'd51;
assign threshold_9[40] = 8'd54;
assign threshold_9[41] = 8'd55;
assign threshold_9[42] = 8'd55;
assign threshold_9[43] = 8'd56;
assign threshold_9[44] = 8'd57;
assign threshold_9[45] = 8'd56;
assign threshold_9[46] = 8'd57;
assign threshold_9[47] = 8'd57;
assign threshold_9[48] = 8'd55;
assign threshold_9[49] = 8'd55;
assign threshold_9[50] = 8'd54;
assign threshold_9[51] = 8'd53;
assign threshold_9[52] = 8'd52;
assign threshold_9[53] = 8'd49;
assign threshold_9[54] = 8'd48;
assign threshold_9[55] = 8'd47;
assign threshold_9[56] = 8'd47;
assign threshold_9[57] = 8'd45;
assign threshold_9[58] = 8'd44;
assign threshold_9[59] = 8'd44;
assign threshold_9[60] = 8'd43;
assign threshold_9[61] = 8'd43;
assign threshold_9[62] = 8'd42;
assign threshold_9[63] = 8'd42;
logic [types::THRESH_BITS-1:0] threshold_10 [64];
assign threshold_10[0] = 8'd58;
assign threshold_10[1] = 8'd58;
assign threshold_10[2] = 8'd57;
assign threshold_10[3] = 8'd55;
assign threshold_10[4] = 8'd53;
assign threshold_10[5] = 8'd51;
assign threshold_10[6] = 8'd47;
assign threshold_10[7] = 8'd44;
assign threshold_10[8] = 8'd40;
assign threshold_10[9] = 8'd35;
assign threshold_10[10] = 8'd31;
assign threshold_10[11] = 8'd26;
assign threshold_10[12] = 8'd21;
assign threshold_10[13] = 8'd15;
assign threshold_10[14] = 8'd11;
assign threshold_10[15] = 8'd5;
assign threshold_10[16] = 8'd0;
assign threshold_10[17] = 8'd5;
assign threshold_10[18] = 8'd9;
assign threshold_10[19] = 8'd14;
assign threshold_10[20] = 8'd18;
assign threshold_10[21] = 8'd22;
assign threshold_10[22] = 8'd25;
assign threshold_10[23] = 8'd29;
assign threshold_10[24] = 8'd31;
assign threshold_10[25] = 8'd34;
assign threshold_10[26] = 8'd36;
assign threshold_10[27] = 8'd38;
assign threshold_10[28] = 8'd40;
assign threshold_10[29] = 8'd41;
assign threshold_10[30] = 8'd41;
assign threshold_10[31] = 8'd41;
assign threshold_10[32] = 8'd42;
assign threshold_10[33] = 8'd42;
assign threshold_10[34] = 8'd41;
assign threshold_10[35] = 8'd41;
assign threshold_10[36] = 8'd40;
assign threshold_10[37] = 8'd38;
assign threshold_10[38] = 8'd37;
assign threshold_10[39] = 8'd34;
assign threshold_10[40] = 8'd31;
assign threshold_10[41] = 8'd29;
assign threshold_10[42] = 8'd26;
assign threshold_10[43] = 8'd22;
assign threshold_10[44] = 8'd18;
assign threshold_10[45] = 8'd14;
assign threshold_10[46] = 8'd10;
assign threshold_10[47] = 8'd5;
assign threshold_10[48] = 8'd0;
assign threshold_10[49] = 8'd5;
assign threshold_10[50] = 8'd10;
assign threshold_10[51] = 8'd15;
assign threshold_10[52] = 8'd20;
assign threshold_10[53] = 8'd26;
assign threshold_10[54] = 8'd30;
assign threshold_10[55] = 8'd36;
assign threshold_10[56] = 8'd39;
assign threshold_10[57] = 8'd44;
assign threshold_10[58] = 8'd47;
assign threshold_10[59] = 8'd50;
assign threshold_10[60] = 8'd54;
assign threshold_10[61] = 8'd55;
assign threshold_10[62] = 8'd56;
assign threshold_10[63] = 8'd58;
logic [types::THRESH_BITS-1:0] threshold_11 [64];
assign threshold_11[0] = 8'd0;
assign threshold_11[1] = 8'd6;
assign threshold_11[2] = 8'd11;
assign threshold_11[3] = 8'd17;
assign threshold_11[4] = 8'd23;
assign threshold_11[5] = 8'd28;
assign threshold_11[6] = 8'd33;
assign threshold_11[7] = 8'd37;
assign threshold_11[8] = 8'd41;
assign threshold_11[9] = 8'd45;
assign threshold_11[10] = 8'd49;
assign threshold_11[11] = 8'd51;
assign threshold_11[12] = 8'd53;
assign threshold_11[13] = 8'd54;
assign threshold_11[14] = 8'd56;
assign threshold_11[15] = 8'd56;
assign threshold_11[16] = 8'd55;
assign threshold_11[17] = 8'd56;
assign threshold_11[18] = 8'd54;
assign threshold_11[19] = 8'd53;
assign threshold_11[20] = 8'd52;
assign threshold_11[21] = 8'd50;
assign threshold_11[22] = 8'd49;
assign threshold_11[23] = 8'd47;
assign threshold_11[24] = 8'd45;
assign threshold_11[25] = 8'd43;
assign threshold_11[26] = 8'd41;
assign threshold_11[27] = 8'd41;
assign threshold_11[28] = 8'd41;
assign threshold_11[29] = 8'd39;
assign threshold_11[30] = 8'd40;
assign threshold_11[31] = 8'd40;
assign threshold_11[32] = 8'd41;
assign threshold_11[33] = 8'd42;
assign threshold_11[34] = 8'd43;
assign threshold_11[35] = 8'd45;
assign threshold_11[36] = 8'd46;
assign threshold_11[37] = 8'd49;
assign threshold_11[38] = 8'd50;
assign threshold_11[39] = 8'd52;
assign threshold_11[40] = 8'd53;
assign threshold_11[41] = 8'd55;
assign threshold_11[42] = 8'd55;
assign threshold_11[43] = 8'd56;
assign threshold_11[44] = 8'd56;
assign threshold_11[45] = 8'd57;
assign threshold_11[46] = 8'd57;
assign threshold_11[47] = 8'd57;
assign threshold_11[48] = 8'd55;
assign threshold_11[49] = 8'd54;
assign threshold_11[50] = 8'd54;
assign threshold_11[51] = 8'd52;
assign threshold_11[52] = 8'd52;
assign threshold_11[53] = 8'd50;
assign threshold_11[54] = 8'd48;
assign threshold_11[55] = 8'd47;
assign threshold_11[56] = 8'd45;
assign threshold_11[57] = 8'd45;
assign threshold_11[58] = 8'd44;
assign threshold_11[59] = 8'd43;
assign threshold_11[60] = 8'd42;
assign threshold_11[61] = 8'd43;
assign threshold_11[62] = 8'd42;
assign threshold_11[63] = 8'd42;

endmodule
